magic
tech sky130A
timestamp 1616337554
<< nwell >>
rect 660 230 2410 660
rect 2050 0 2410 230
<< nmos >>
rect 810 30 860 150
rect 1010 30 1060 150
rect 1120 30 1170 150
rect 1470 30 1520 150
rect 1690 30 1740 150
rect 1800 30 1850 150
rect 1280 -220 1330 -100
rect 1480 -220 1530 -100
rect 1590 -220 1640 -100
rect 1790 -220 1840 -100
rect 1900 -220 1950 -100
rect 2200 -220 2250 -100
<< pmos >>
rect 810 500 860 620
rect 1060 500 1110 620
rect 1170 500 1220 620
rect 1370 500 1420 620
rect 1480 500 1530 620
rect 1740 500 1790 620
rect 2000 500 2050 620
rect 2200 500 2250 620
rect 810 270 860 390
rect 1010 270 1060 390
rect 1270 270 1320 390
rect 1380 270 1430 390
rect 1580 270 1630 390
rect 1690 270 1740 390
rect 2000 270 2050 390
rect 2200 270 2250 390
rect 2130 40 2180 160
<< ndiff >>
rect 750 130 810 150
rect 750 50 770 130
rect 790 50 810 130
rect 750 30 810 50
rect 860 130 920 150
rect 860 50 880 130
rect 900 50 920 130
rect 860 30 920 50
rect 950 130 1010 150
rect 950 50 970 130
rect 990 50 1010 130
rect 950 30 1010 50
rect 1060 130 1120 150
rect 1060 50 1080 130
rect 1100 50 1120 130
rect 1060 30 1120 50
rect 1170 130 1230 150
rect 1170 50 1190 130
rect 1210 50 1230 130
rect 1170 30 1230 50
rect 1410 130 1470 150
rect 1410 50 1430 130
rect 1450 50 1470 130
rect 1410 30 1470 50
rect 1520 130 1580 150
rect 1520 50 1540 130
rect 1560 50 1580 130
rect 1520 30 1580 50
rect 1630 130 1690 150
rect 1630 50 1650 130
rect 1670 50 1690 130
rect 1630 30 1690 50
rect 1740 130 1800 150
rect 1740 50 1760 130
rect 1780 50 1800 130
rect 1740 30 1800 50
rect 1850 130 1910 150
rect 1850 50 1870 130
rect 1890 50 1910 130
rect 1850 30 1910 50
rect 1220 -120 1280 -100
rect 1220 -200 1240 -120
rect 1260 -200 1280 -120
rect 1220 -220 1280 -200
rect 1330 -120 1390 -100
rect 1330 -200 1350 -120
rect 1370 -200 1390 -120
rect 1330 -220 1390 -200
rect 1420 -120 1480 -100
rect 1420 -200 1440 -120
rect 1460 -200 1480 -120
rect 1420 -220 1480 -200
rect 1530 -120 1590 -100
rect 1530 -200 1550 -120
rect 1570 -200 1590 -120
rect 1530 -220 1590 -200
rect 1640 -120 1700 -100
rect 1640 -200 1660 -120
rect 1680 -200 1700 -120
rect 1640 -220 1700 -200
rect 1730 -120 1790 -100
rect 1730 -200 1750 -120
rect 1770 -200 1790 -120
rect 1730 -220 1790 -200
rect 1840 -120 1900 -100
rect 1840 -200 1860 -120
rect 1880 -200 1900 -120
rect 1840 -220 1900 -200
rect 1950 -120 2010 -100
rect 1950 -200 1970 -120
rect 1990 -200 2010 -120
rect 1950 -220 2010 -200
rect 2140 -120 2200 -100
rect 2140 -200 2160 -120
rect 2180 -200 2200 -120
rect 2140 -220 2200 -200
rect 2250 -120 2310 -100
rect 2250 -200 2270 -120
rect 2290 -200 2310 -120
rect 2250 -220 2310 -200
<< pdiff >>
rect 750 600 810 620
rect 750 520 770 600
rect 790 520 810 600
rect 750 500 810 520
rect 860 600 920 620
rect 860 520 880 600
rect 900 520 920 600
rect 860 500 920 520
rect 1000 600 1060 620
rect 1000 520 1020 600
rect 1040 520 1060 600
rect 1000 500 1060 520
rect 1110 600 1170 620
rect 1110 520 1130 600
rect 1150 520 1170 600
rect 1110 500 1170 520
rect 1220 600 1280 620
rect 1220 520 1240 600
rect 1260 520 1280 600
rect 1220 500 1280 520
rect 1310 600 1370 620
rect 1310 520 1330 600
rect 1350 520 1370 600
rect 1310 500 1370 520
rect 1420 600 1480 620
rect 1420 520 1440 600
rect 1460 520 1480 600
rect 1420 500 1480 520
rect 1530 600 1590 620
rect 1530 520 1550 600
rect 1570 520 1590 600
rect 1530 500 1590 520
rect 1680 600 1740 620
rect 1680 520 1700 600
rect 1720 520 1740 600
rect 1680 500 1740 520
rect 1790 600 1850 620
rect 1790 520 1810 600
rect 1830 520 1850 600
rect 1790 500 1850 520
rect 1940 600 2000 620
rect 1940 520 1960 600
rect 1980 520 2000 600
rect 1940 500 2000 520
rect 2050 600 2110 620
rect 2050 520 2070 600
rect 2090 520 2110 600
rect 2050 500 2110 520
rect 2140 600 2200 620
rect 2140 520 2160 600
rect 2180 520 2200 600
rect 2140 500 2200 520
rect 2250 600 2310 620
rect 2250 520 2270 600
rect 2290 520 2310 600
rect 2250 500 2310 520
rect 750 370 810 390
rect 750 290 770 370
rect 790 290 810 370
rect 750 270 810 290
rect 860 370 920 390
rect 860 290 880 370
rect 900 290 920 370
rect 860 270 920 290
rect 950 370 1010 390
rect 950 290 970 370
rect 990 290 1010 370
rect 950 270 1010 290
rect 1060 370 1120 390
rect 1060 290 1080 370
rect 1100 290 1120 370
rect 1060 270 1120 290
rect 1210 370 1270 390
rect 1210 290 1230 370
rect 1250 290 1270 370
rect 1210 270 1270 290
rect 1320 370 1380 390
rect 1320 290 1340 370
rect 1360 290 1380 370
rect 1320 270 1380 290
rect 1430 370 1490 390
rect 1430 290 1450 370
rect 1470 290 1490 370
rect 1430 270 1490 290
rect 1520 370 1580 390
rect 1520 290 1540 370
rect 1560 290 1580 370
rect 1520 270 1580 290
rect 1630 370 1690 390
rect 1630 290 1650 370
rect 1670 290 1690 370
rect 1630 270 1690 290
rect 1740 370 1800 390
rect 1740 290 1760 370
rect 1780 290 1800 370
rect 1740 270 1800 290
rect 1940 370 2000 390
rect 1940 290 1960 370
rect 1980 290 2000 370
rect 1940 270 2000 290
rect 2050 370 2110 390
rect 2050 290 2070 370
rect 2090 290 2110 370
rect 2050 270 2110 290
rect 2140 370 2200 390
rect 2140 290 2160 370
rect 2180 290 2200 370
rect 2140 270 2200 290
rect 2250 370 2310 390
rect 2250 290 2270 370
rect 2290 290 2310 370
rect 2250 270 2310 290
rect 2070 140 2130 160
rect 2070 60 2090 140
rect 2110 60 2130 140
rect 2070 40 2130 60
rect 2180 140 2240 160
rect 2180 60 2200 140
rect 2220 60 2240 140
rect 2180 40 2240 60
<< ndiffc >>
rect 770 50 790 130
rect 880 50 900 130
rect 970 50 990 130
rect 1080 50 1100 130
rect 1190 50 1210 130
rect 1430 50 1450 130
rect 1540 50 1560 130
rect 1650 50 1670 130
rect 1760 50 1780 130
rect 1870 50 1890 130
rect 1240 -200 1260 -120
rect 1350 -200 1370 -120
rect 1440 -200 1460 -120
rect 1550 -200 1570 -120
rect 1660 -200 1680 -120
rect 1750 -200 1770 -120
rect 1860 -200 1880 -120
rect 1970 -200 1990 -120
rect 2160 -200 2180 -120
rect 2270 -200 2290 -120
<< pdiffc >>
rect 770 520 790 600
rect 880 520 900 600
rect 1020 520 1040 600
rect 1130 520 1150 600
rect 1240 520 1260 600
rect 1330 520 1350 600
rect 1440 520 1460 600
rect 1550 520 1570 600
rect 1700 520 1720 600
rect 1810 520 1830 600
rect 1960 520 1980 600
rect 2070 520 2090 600
rect 2160 520 2180 600
rect 2270 520 2290 600
rect 770 290 790 370
rect 880 290 900 370
rect 970 290 990 370
rect 1080 290 1100 370
rect 1230 290 1250 370
rect 1340 290 1360 370
rect 1450 290 1470 370
rect 1540 290 1560 370
rect 1650 290 1670 370
rect 1760 290 1780 370
rect 1960 290 1980 370
rect 2070 290 2090 370
rect 2160 290 2180 370
rect 2270 290 2290 370
rect 2090 60 2110 140
rect 2200 60 2220 140
<< psubdiff >>
rect 690 130 750 150
rect 690 50 710 130
rect 730 50 750 130
rect 690 30 750 50
rect 1230 130 1290 150
rect 1230 50 1250 130
rect 1270 50 1290 130
rect 1230 30 1290 50
rect 1350 130 1410 150
rect 1350 50 1370 130
rect 1390 50 1410 130
rect 1350 30 1410 50
rect 1160 -120 1220 -100
rect 1160 -200 1180 -120
rect 1200 -200 1220 -120
rect 1160 -220 1220 -200
rect 2310 -120 2370 -100
rect 2310 -200 2330 -120
rect 2350 -200 2370 -120
rect 2310 -220 2370 -200
<< nsubdiff >>
rect 690 600 750 620
rect 690 520 710 600
rect 730 520 750 600
rect 690 500 750 520
rect 1620 600 1680 620
rect 1620 520 1640 600
rect 1660 520 1680 600
rect 1620 500 1680 520
rect 1880 600 1940 620
rect 1880 520 1900 600
rect 1920 520 1940 600
rect 1880 500 1940 520
rect 2310 600 2370 620
rect 2310 520 2330 600
rect 2350 520 2370 600
rect 2310 500 2370 520
rect 690 370 750 390
rect 690 290 710 370
rect 730 290 750 370
rect 690 270 750 290
rect 1120 370 1180 390
rect 1120 290 1140 370
rect 1160 290 1180 370
rect 1120 270 1180 290
rect 1880 370 1940 390
rect 1880 290 1900 370
rect 1920 290 1940 370
rect 1880 270 1940 290
rect 2310 370 2370 390
rect 2310 290 2330 370
rect 2350 290 2370 370
rect 2310 270 2370 290
rect 2240 140 2300 160
rect 2240 60 2260 140
rect 2280 60 2300 140
rect 2240 40 2300 60
<< psubdiffcont >>
rect 710 50 730 130
rect 1250 50 1270 130
rect 1370 50 1390 130
rect 1180 -200 1200 -120
rect 2330 -200 2350 -120
<< nsubdiffcont >>
rect 710 520 730 600
rect 1640 520 1660 600
rect 1900 520 1920 600
rect 2330 520 2350 600
rect 710 290 730 370
rect 1140 290 1160 370
rect 1900 290 1920 370
rect 2330 290 2350 370
rect 2260 60 2280 140
<< poly >>
rect 1560 700 1600 710
rect 1560 690 1570 700
rect 930 680 1570 690
rect 1590 690 1600 700
rect 1590 680 2320 690
rect 930 660 940 680
rect 960 670 2290 680
rect 960 660 970 670
rect 930 650 970 660
rect 810 620 860 640
rect 1060 620 1110 670
rect 1180 640 1210 670
rect 1380 640 1410 670
rect 1490 640 1520 670
rect 1750 640 1780 670
rect 2280 660 2290 670
rect 2310 660 2320 680
rect 2280 650 2320 660
rect 1170 620 1220 640
rect 1370 620 1420 640
rect 1480 620 1530 640
rect 1740 620 1790 640
rect 2000 620 2050 640
rect 2200 620 2250 640
rect 810 490 860 500
rect 700 480 860 490
rect 1060 480 1110 500
rect 1170 480 1220 500
rect 1370 480 1420 500
rect 1480 480 1530 500
rect 1740 480 1790 500
rect 700 460 710 480
rect 730 470 860 480
rect 730 460 740 470
rect 700 450 740 460
rect 1490 450 1520 480
rect 1010 430 1740 450
rect 810 390 860 410
rect 1010 390 1060 430
rect 1270 390 1320 430
rect 1380 390 1430 430
rect 1580 390 1630 430
rect 1690 390 1740 430
rect 1890 440 1930 450
rect 2000 440 2050 500
rect 2200 480 2250 500
rect 1890 420 1900 440
rect 1920 420 2050 440
rect 1890 410 1930 420
rect 2000 390 2050 420
rect 2200 390 2250 410
rect 810 250 860 270
rect 1010 250 1060 270
rect 1270 250 1320 270
rect 1380 250 1430 270
rect 1580 250 1630 270
rect 1690 250 1740 270
rect 2000 250 2050 270
rect 2200 250 2250 270
rect 700 240 860 250
rect 700 220 710 240
rect 730 230 860 240
rect 730 220 740 230
rect 700 210 740 220
rect 2130 210 2250 220
rect 960 200 1000 210
rect 960 180 970 200
rect 990 190 1000 200
rect 1550 200 1590 210
rect 1550 190 1560 200
rect 990 180 1060 190
rect 960 170 1060 180
rect 1470 180 1560 190
rect 1580 180 1590 200
rect 1470 170 1590 180
rect 1620 200 1660 210
rect 2130 200 2220 210
rect 1620 180 1630 200
rect 1650 180 1740 200
rect 1620 170 1660 180
rect 810 150 860 170
rect 1010 150 1060 170
rect 1120 150 1170 170
rect 1470 150 1520 170
rect 1690 150 1740 180
rect 1800 150 1850 170
rect 2130 160 2180 200
rect 2210 190 2220 200
rect 2240 190 2250 210
rect 2210 180 2250 190
rect 810 10 860 30
rect 700 0 860 10
rect 700 -20 710 0
rect 730 -10 860 0
rect 1010 10 1060 30
rect 1120 10 1170 30
rect 1470 10 1520 30
rect 1010 -10 1170 10
rect 730 -20 740 -10
rect 700 -30 740 -20
rect 1690 -60 1740 30
rect 1800 10 1850 30
rect 2130 20 2180 40
rect 1910 0 1950 10
rect 1910 -20 1920 0
rect 1940 -10 1950 0
rect 2240 0 2280 10
rect 2240 -10 2250 0
rect 1940 -20 2250 -10
rect 2270 -20 2280 0
rect 1910 -30 2280 -20
rect 1480 -70 2120 -60
rect 1480 -80 2090 -70
rect 1280 -100 1330 -80
rect 1480 -100 1530 -80
rect 1590 -100 1640 -80
rect 1790 -100 1840 -80
rect 1900 -100 1950 -80
rect 2080 -90 2090 -80
rect 2110 -90 2120 -70
rect 2080 -100 2120 -90
rect 2200 -100 2250 -80
rect 1280 -240 1330 -220
rect 1480 -240 1530 -220
rect 1590 -240 1640 -220
rect 1790 -240 1840 -220
rect 1900 -240 1950 -220
rect 2200 -240 2250 -220
rect 1170 -250 1330 -240
rect 1170 -270 1180 -250
rect 1200 -260 1330 -250
rect 2200 -250 2360 -240
rect 2200 -260 2330 -250
rect 1200 -270 1210 -260
rect 1170 -280 1210 -270
rect 2320 -270 2330 -260
rect 2350 -270 2360 -250
rect 2320 -280 2360 -270
<< polycont >>
rect 1570 680 1590 700
rect 940 660 960 680
rect 2290 660 2310 680
rect 710 460 730 480
rect 1900 420 1920 440
rect 710 220 730 240
rect 970 180 990 200
rect 1560 180 1580 200
rect 1630 180 1650 200
rect 2220 190 2240 210
rect 710 -20 730 0
rect 1920 -20 1940 0
rect 2250 -20 2270 0
rect 2090 -90 2110 -70
rect 1180 -270 1200 -250
rect 2330 -270 2350 -250
<< locali >>
rect 1560 700 1600 710
rect 660 680 970 690
rect 660 660 940 680
rect 960 660 970 680
rect 1560 680 1570 700
rect 1590 680 1600 700
rect 1560 670 1600 680
rect 2280 680 2410 690
rect 660 650 970 660
rect 1140 640 1450 660
rect 1140 610 1160 640
rect 1430 610 1450 640
rect 1560 610 1580 670
rect 2280 660 2290 680
rect 2310 660 2410 680
rect 2280 650 2320 660
rect 700 600 800 610
rect 700 520 710 600
rect 730 520 770 600
rect 790 520 800 600
rect 700 510 800 520
rect 870 600 1050 610
rect 870 520 880 600
rect 900 590 1020 600
rect 900 520 910 590
rect 870 510 910 520
rect 1010 520 1020 590
rect 1040 520 1050 600
rect 1010 510 1050 520
rect 1120 600 1160 610
rect 1120 520 1130 600
rect 1150 520 1160 600
rect 1120 510 1160 520
rect 1230 600 1270 610
rect 1230 520 1240 600
rect 1260 520 1270 600
rect 1230 510 1270 520
rect 700 490 720 510
rect 700 480 740 490
rect 700 460 710 480
rect 730 460 740 480
rect 1030 480 1050 510
rect 1250 480 1270 510
rect 1320 600 1360 610
rect 1320 520 1330 600
rect 1350 520 1360 600
rect 1320 510 1360 520
rect 1430 600 1470 610
rect 1430 520 1440 600
rect 1460 520 1470 600
rect 1430 510 1470 520
rect 1540 600 1580 610
rect 1540 520 1550 600
rect 1570 520 1580 600
rect 1540 510 1580 520
rect 1630 600 1730 610
rect 1630 520 1640 600
rect 1660 520 1700 600
rect 1720 520 1730 600
rect 1630 510 1730 520
rect 1800 600 1840 610
rect 1800 520 1810 600
rect 1830 520 1840 600
rect 1800 510 1840 520
rect 1890 600 1990 610
rect 1890 520 1900 600
rect 1920 520 1960 600
rect 1980 520 1990 600
rect 1890 510 1990 520
rect 2060 600 2190 610
rect 2060 520 2070 600
rect 2090 590 2160 600
rect 2090 520 2100 590
rect 2060 510 2100 520
rect 2150 520 2160 590
rect 2180 520 2190 600
rect 2150 510 2190 520
rect 2260 600 2360 610
rect 2260 520 2270 600
rect 2290 520 2330 600
rect 2350 520 2360 600
rect 2260 510 2360 520
rect 1320 480 1340 510
rect 1540 480 1560 510
rect 1030 460 1560 480
rect 700 450 740 460
rect 1350 410 1660 430
rect 1350 380 1370 410
rect 1640 380 1660 410
rect 700 370 800 380
rect 700 290 710 370
rect 730 290 770 370
rect 790 290 800 370
rect 700 280 800 290
rect 870 370 1000 380
rect 870 290 880 370
rect 900 360 970 370
rect 900 290 910 360
rect 870 280 910 290
rect 960 290 970 360
rect 990 290 1000 370
rect 960 280 1000 290
rect 1070 370 1170 380
rect 1070 290 1080 370
rect 1100 290 1140 370
rect 1160 290 1170 370
rect 1070 280 1170 290
rect 1220 370 1260 380
rect 1220 290 1230 370
rect 1250 290 1260 370
rect 1220 280 1260 290
rect 1330 370 1370 380
rect 1330 290 1340 370
rect 1360 290 1370 370
rect 1330 280 1370 290
rect 1440 370 1480 380
rect 1440 290 1450 370
rect 1470 290 1480 370
rect 1440 280 1480 290
rect 700 250 720 280
rect 700 240 740 250
rect 700 220 710 240
rect 730 220 740 240
rect 700 210 740 220
rect 960 210 980 280
rect 1240 250 1260 280
rect 1460 250 1480 280
rect 1530 370 1570 380
rect 1530 290 1540 370
rect 1560 290 1570 370
rect 1530 280 1570 290
rect 1640 370 1680 380
rect 1640 290 1650 370
rect 1670 290 1680 370
rect 1640 280 1680 290
rect 1750 370 1790 380
rect 1750 290 1760 370
rect 1780 290 1790 370
rect 1750 280 1790 290
rect 1530 250 1550 280
rect 1750 250 1770 280
rect 1240 230 1770 250
rect 1550 210 1570 230
rect 960 200 1000 210
rect 960 180 970 200
rect 990 180 1000 200
rect 960 170 1000 180
rect 1550 200 1590 210
rect 1550 180 1560 200
rect 1580 180 1590 200
rect 1550 170 1590 180
rect 1620 200 1660 210
rect 1810 200 1830 510
rect 1890 440 1930 450
rect 1890 420 1900 440
rect 1920 420 1930 440
rect 1890 410 1930 420
rect 1900 380 1920 410
rect 2060 380 2080 510
rect 1890 370 1990 380
rect 1890 300 1900 370
rect 1620 180 1630 200
rect 1650 180 1830 200
rect 1860 290 1900 300
rect 1920 290 1960 370
rect 1980 290 1990 370
rect 1860 280 1990 290
rect 2060 370 2190 380
rect 2060 290 2070 370
rect 2090 360 2160 370
rect 2090 290 2100 360
rect 2060 280 2100 290
rect 2150 290 2160 360
rect 2180 290 2190 370
rect 2150 280 2190 290
rect 2260 370 2360 380
rect 2260 290 2270 370
rect 2290 290 2330 370
rect 2350 290 2360 370
rect 2260 280 2360 290
rect 1620 170 1660 180
rect 960 140 980 170
rect 1550 140 1570 170
rect 700 130 800 140
rect 700 50 710 130
rect 730 50 770 130
rect 790 50 800 130
rect 700 40 800 50
rect 870 130 1000 140
rect 870 50 880 130
rect 900 120 970 130
rect 900 50 910 120
rect 870 40 910 50
rect 960 50 970 120
rect 990 50 1000 130
rect 960 40 1000 50
rect 1070 130 1110 140
rect 1070 50 1080 130
rect 1100 50 1110 130
rect 1070 40 1110 50
rect 1180 130 1280 140
rect 1180 50 1190 130
rect 1210 50 1250 130
rect 1270 50 1280 130
rect 1180 40 1280 50
rect 1360 130 1460 140
rect 1360 50 1370 130
rect 1390 50 1430 130
rect 1450 50 1460 130
rect 1360 40 1460 50
rect 1530 130 1570 140
rect 1530 50 1540 130
rect 1560 50 1570 130
rect 1530 40 1570 50
rect 1640 140 1660 170
rect 1860 140 1880 280
rect 2080 150 2100 280
rect 2210 210 2250 220
rect 2210 190 2220 210
rect 2240 190 2250 210
rect 2210 180 2250 190
rect 2210 150 2230 180
rect 2080 140 2120 150
rect 1640 130 1680 140
rect 1640 50 1650 130
rect 1670 50 1680 130
rect 1640 40 1680 50
rect 1750 130 1790 140
rect 1750 50 1760 130
rect 1780 50 1790 130
rect 1750 40 1790 50
rect 1860 130 1900 140
rect 1860 50 1870 130
rect 1890 50 1900 130
rect 2080 60 2090 140
rect 2110 60 2120 140
rect 2080 50 2120 60
rect 2190 140 2410 150
rect 2190 60 2200 140
rect 2220 60 2260 140
rect 2280 120 2410 140
rect 2280 60 2290 120
rect 2190 50 2290 60
rect 1860 40 1900 50
rect 700 10 720 40
rect 1090 10 1110 40
rect 1360 10 1380 40
rect 700 0 740 10
rect 700 -20 710 0
rect 730 -20 740 0
rect 1090 -10 1380 10
rect 1540 10 1570 40
rect 2190 10 2210 50
rect 1540 0 1950 10
rect 1540 -20 1920 0
rect 1940 -20 1950 0
rect 700 -30 740 -20
rect 1910 -30 1950 -20
rect 1980 -10 2210 10
rect 2240 0 2410 10
rect 1980 -110 2000 -10
rect 2240 -20 2250 0
rect 2270 -20 2410 0
rect 2240 -30 2280 -20
rect 2080 -70 2410 -60
rect 2080 -90 2090 -70
rect 2110 -90 2410 -70
rect 2080 -100 2120 -90
rect 1170 -120 1270 -110
rect 1170 -200 1180 -120
rect 1200 -200 1240 -120
rect 1260 -200 1270 -120
rect 1170 -210 1270 -200
rect 1340 -120 1470 -110
rect 1340 -200 1350 -120
rect 1370 -130 1440 -120
rect 1370 -200 1380 -130
rect 1340 -210 1380 -200
rect 1430 -200 1440 -130
rect 1460 -200 1470 -120
rect 1430 -210 1470 -200
rect 1540 -120 1580 -110
rect 1540 -200 1550 -120
rect 1570 -200 1580 -120
rect 1540 -210 1580 -200
rect 1650 -120 1690 -110
rect 1650 -200 1660 -120
rect 1680 -200 1690 -120
rect 1650 -210 1690 -200
rect 1170 -240 1190 -210
rect 1450 -240 1470 -210
rect 1670 -240 1690 -210
rect 1740 -120 1780 -110
rect 1740 -200 1750 -120
rect 1770 -200 1780 -120
rect 1740 -210 1780 -200
rect 1850 -120 1890 -110
rect 1850 -200 1860 -120
rect 1880 -200 1890 -120
rect 1850 -210 1890 -200
rect 1960 -120 2000 -110
rect 1960 -200 1970 -120
rect 1990 -190 2000 -120
rect 2150 -120 2190 -110
rect 2150 -190 2160 -120
rect 1990 -200 2160 -190
rect 2180 -200 2190 -120
rect 1960 -210 2190 -200
rect 2260 -120 2360 -110
rect 2260 -200 2270 -120
rect 2290 -200 2330 -120
rect 2350 -200 2360 -120
rect 2260 -210 2360 -200
rect 1740 -240 1760 -210
rect 1960 -240 1980 -210
rect 2340 -240 2360 -210
rect 1170 -250 1210 -240
rect 1170 -270 1180 -250
rect 1200 -270 1210 -250
rect 1450 -260 1980 -240
rect 2320 -250 2360 -240
rect 1170 -280 1210 -270
rect 2320 -270 2330 -250
rect 2350 -270 2360 -250
rect 2320 -280 2360 -270
<< viali >>
rect 710 520 730 600
rect 770 520 790 600
rect 1130 520 1150 600
rect 1440 520 1460 600
rect 1640 520 1660 600
rect 1700 520 1720 600
rect 1900 520 1920 600
rect 1960 520 1980 600
rect 2270 520 2290 600
rect 2330 520 2350 600
rect 710 290 730 370
rect 770 290 790 370
rect 1080 290 1100 370
rect 1140 290 1160 370
rect 1340 290 1360 370
rect 1650 290 1670 370
rect 2270 290 2290 370
rect 2330 290 2350 370
rect 710 50 730 130
rect 770 50 790 130
rect 1190 50 1210 130
rect 1250 50 1270 130
rect 1760 50 1780 130
rect 1180 -200 1200 -120
rect 1240 -200 1260 -120
rect 1550 -200 1570 -120
rect 1860 -200 1880 -120
rect 2270 -200 2290 -120
rect 2330 -200 2350 -120
<< metal1 >>
rect 1560 610 1580 650
rect 660 600 2410 610
rect 660 520 710 600
rect 730 520 770 600
rect 790 520 1130 600
rect 1150 520 1440 600
rect 1460 520 1640 600
rect 1660 520 1700 600
rect 1720 520 1900 600
rect 1920 520 1960 600
rect 1980 520 2270 600
rect 2290 520 2330 600
rect 2350 520 2410 600
rect 660 370 2410 520
rect 660 290 710 370
rect 730 290 770 370
rect 790 290 1080 370
rect 1100 290 1140 370
rect 1160 290 1340 370
rect 1360 290 1650 370
rect 1670 290 2270 370
rect 2290 290 2330 370
rect 2350 290 2410 370
rect 660 280 2410 290
rect 660 130 2410 160
rect 660 50 710 130
rect 730 50 770 130
rect 790 50 1190 130
rect 1210 50 1250 130
rect 1270 50 1760 130
rect 1780 50 2410 130
rect 660 -120 2410 50
rect 660 -200 1180 -120
rect 1200 -200 1240 -120
rect 1260 -200 1550 -120
rect 1570 -200 1860 -120
rect 1880 -200 2270 -120
rect 2290 -200 2330 -120
rect 2350 -200 2410 -120
rect 660 -210 2410 -200
<< labels >>
rlabel metal1 660 -20 660 -20 7 VN
rlabel metal1 660 440 660 440 7 VP
rlabel locali 660 670 660 670 7 Vb
rlabel locali 2410 130 2410 130 3 Vcp
rlabel locali 2410 0 2410 0 3 Vcn
rlabel locali 2410 -70 2410 -70 3 Vbn
<< end >>
