* SPICE3 file created from Amplifier.ext - technology: sky130A


* Top level circuit Amplifier

X0 VP Vbp a_3170_380# VP sky130_fd_pr__pfet_01v8 ad=2.4e+13p pd=1e+08u as=1.2e+13p ps=5e+07u w=1.2e+07u l=500000u
X1 Vout Vcp a_4530_380# VP sky130_fd_pr__pfet_01v8 ad=6e+12p pd=2.5e+07u as=6e+12p ps=2.5e+07u w=1.2e+07u l=500000u
X2 VN VN Vout VN sky130_fd_pr__nfet_01v8 ad=1.8e+13p pd=7.5e+07u as=6e+12p ps=2.5e+07u w=1.2e+07u l=500000u
X3 VP a_3930_n2320# a_4130_380# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6e+12p ps=2.5e+07u w=1.2e+07u l=500000u
X4 a_3930_n2320# VN VN VN sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.5e+07u as=0p ps=0u w=1.2e+07u l=500000u
X5 VP VP Vout VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X6 a_3930_n2320# VP VP VP sky130_fd_pr__pfet_01v8 ad=6e+12p pd=2.5e+07u as=0p ps=0u w=1.2e+07u l=500000u
X7 a_4530_380# a_3930_n2320# VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X8 a_3170_380# V2 a_3010_n2320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=6e+12p ps=2.5e+07u w=1.2e+07u l=500000u
X9 a_3410_n2320# Vcn a_3930_n2320# VN sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.5e+07u as=0p ps=0u w=1.2e+07u l=500000u
X10 a_4130_380# Vcp a_3930_n2320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X11 a_3410_n2320# V1 a_3170_380# VP sky130_fd_pr__pfet_01v8 ad=6e+12p pd=2.5e+07u as=0p ps=0u w=1.2e+07u l=500000u
X12 VN Vbn a_3410_n2320# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
X13 a_3010_n2320# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=6e+12p pd=2.5e+07u as=0p ps=0u w=1.2e+07u l=500000u
X14 Vout Vcn a_3010_n2320# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.2e+07u l=500000u
.end

