magic
tech sky130A
timestamp 1618004850
<< nwell >>
rect 1435 155 2585 1410
rect 1435 -1180 1775 155
<< nmos >>
rect 1915 -1160 1965 40
rect 2015 -1160 2065 40
rect 2115 -1160 2165 40
rect 2215 -1160 2265 40
rect 2315 -1160 2365 40
rect 2415 -1160 2465 40
<< pmos >>
rect 1635 190 1685 1390
rect 1915 190 1965 1390
rect 2015 190 2065 1390
rect 2115 190 2165 1390
rect 2215 190 2265 1390
rect 2315 190 2365 1390
rect 2415 190 2465 1390
rect 1555 -1160 1605 40
rect 1655 -1160 1705 40
<< ndiff >>
rect 1865 25 1915 40
rect 1865 -1145 1880 25
rect 1900 -1145 1915 25
rect 1865 -1160 1915 -1145
rect 1965 25 2015 40
rect 1965 -1145 1980 25
rect 2000 -1145 2015 25
rect 1965 -1160 2015 -1145
rect 2065 25 2115 40
rect 2065 -1145 2080 25
rect 2100 -1145 2115 25
rect 2065 -1160 2115 -1145
rect 2165 25 2215 40
rect 2165 -1145 2180 25
rect 2200 -1145 2215 25
rect 2165 -1160 2215 -1145
rect 2265 25 2315 40
rect 2265 -1145 2280 25
rect 2300 -1145 2315 25
rect 2265 -1160 2315 -1145
rect 2365 25 2415 40
rect 2365 -1145 2380 25
rect 2400 -1145 2415 25
rect 2365 -1160 2415 -1145
rect 2465 25 2515 40
rect 2465 -1145 2480 25
rect 2500 -1145 2515 25
rect 2465 -1160 2515 -1145
<< pdiff >>
rect 1585 1375 1635 1390
rect 1585 205 1600 1375
rect 1620 205 1635 1375
rect 1585 190 1635 205
rect 1685 1375 1735 1390
rect 1685 205 1700 1375
rect 1720 205 1735 1375
rect 1685 190 1735 205
rect 1865 1375 1915 1390
rect 1865 205 1880 1375
rect 1900 205 1915 1375
rect 1865 190 1915 205
rect 1965 1375 2015 1390
rect 1965 205 1980 1375
rect 2000 205 2015 1375
rect 1965 190 2015 205
rect 2065 1375 2115 1390
rect 2065 205 2080 1375
rect 2100 205 2115 1375
rect 2065 190 2115 205
rect 2165 1375 2215 1390
rect 2165 205 2180 1375
rect 2200 205 2215 1375
rect 2165 190 2215 205
rect 2265 1370 2315 1390
rect 2265 210 2280 1370
rect 2300 210 2315 1370
rect 2265 190 2315 210
rect 2365 1375 2415 1390
rect 2365 205 2380 1375
rect 2400 205 2415 1375
rect 2365 190 2415 205
rect 2465 1375 2515 1390
rect 2465 205 2480 1375
rect 2500 205 2515 1375
rect 2465 190 2515 205
rect 1505 25 1555 40
rect 1505 -1145 1520 25
rect 1540 -1145 1555 25
rect 1505 -1160 1555 -1145
rect 1605 25 1655 40
rect 1605 -1145 1620 25
rect 1640 -1145 1655 25
rect 1605 -1160 1655 -1145
rect 1705 25 1755 40
rect 1705 -1145 1720 25
rect 1740 -1145 1755 25
rect 1705 -1160 1755 -1145
<< ndiffc >>
rect 1880 -1145 1900 25
rect 1980 -1145 2000 25
rect 2080 -1145 2100 25
rect 2180 -1145 2200 25
rect 2280 -1145 2300 25
rect 2380 -1145 2400 25
rect 2480 -1145 2500 25
<< pdiffc >>
rect 1600 205 1620 1375
rect 1700 205 1720 1375
rect 1880 205 1900 1375
rect 1980 205 2000 1375
rect 2080 205 2100 1375
rect 2180 205 2200 1375
rect 2280 210 2300 1370
rect 2380 205 2400 1375
rect 2480 205 2500 1375
rect 1520 -1145 1540 25
rect 1620 -1145 1640 25
rect 1720 -1145 1740 25
<< psubdiff >>
rect 1815 25 1865 40
rect 1815 -1145 1830 25
rect 1850 -1145 1865 25
rect 1815 -1160 1865 -1145
rect 2515 25 2565 40
rect 2515 -1145 2530 25
rect 2550 -1145 2565 25
rect 2515 -1160 2565 -1145
<< nsubdiff >>
rect 1735 1375 1785 1390
rect 1735 205 1750 1375
rect 1770 205 1785 1375
rect 1735 190 1785 205
rect 1815 1375 1865 1390
rect 1815 205 1830 1375
rect 1850 205 1865 1375
rect 1815 190 1865 205
rect 2515 1375 2565 1390
rect 2515 205 2530 1375
rect 2550 205 2565 1375
rect 2515 190 2565 205
<< psubdiffcont >>
rect 1830 -1145 1850 25
rect 2530 -1145 2550 25
<< nsubdiffcont >>
rect 1750 205 1770 1375
rect 1830 205 1850 1375
rect 2530 205 2550 1375
<< poly >>
rect 2170 1480 2210 1490
rect 2170 1460 2180 1480
rect 2200 1460 2210 1480
rect 2170 1450 2210 1460
rect 1870 1435 1910 1445
rect 1530 1410 1685 1420
rect 1530 1390 1540 1410
rect 1560 1405 1685 1410
rect 1870 1415 1880 1435
rect 1900 1420 1910 1435
rect 2015 1430 2365 1450
rect 1900 1415 1965 1420
rect 1870 1405 1965 1415
rect 1560 1390 1570 1405
rect 1635 1390 1685 1405
rect 1915 1390 1965 1405
rect 2015 1390 2065 1430
rect 2115 1390 2165 1405
rect 2215 1390 2265 1405
rect 2315 1390 2365 1430
rect 2470 1435 2510 1445
rect 2470 1420 2480 1435
rect 2415 1415 2480 1420
rect 2500 1415 2510 1435
rect 2415 1405 2510 1415
rect 2415 1390 2465 1405
rect 1530 1380 1570 1390
rect 1635 175 1685 190
rect 1915 175 1965 190
rect 2015 175 2065 190
rect 2115 175 2165 190
rect 2215 175 2265 190
rect 2315 175 2365 190
rect 2415 175 2465 190
rect 2115 165 2265 175
rect 2115 160 2180 165
rect 1550 150 1590 160
rect 1550 130 1560 150
rect 1580 135 1590 150
rect 2170 145 2180 160
rect 2200 160 2265 165
rect 2200 145 2210 160
rect 2170 135 2210 145
rect 1580 130 2130 135
rect 1550 120 2130 130
rect 1490 85 2065 95
rect 1490 65 1500 85
rect 1520 80 2065 85
rect 1520 65 1530 80
rect 1490 55 1530 65
rect 1555 40 1605 55
rect 1655 40 1705 55
rect 1915 40 1965 55
rect 2015 40 2065 80
rect 2115 75 2130 120
rect 2115 55 2265 75
rect 2115 40 2165 55
rect 2215 40 2265 55
rect 2315 40 2365 55
rect 2415 40 2465 55
rect 1450 -1160 1490 -1150
rect 1450 -1180 1460 -1160
rect 1480 -1175 1490 -1160
rect 1555 -1175 1605 -1160
rect 1480 -1180 1605 -1175
rect 1450 -1190 1605 -1180
rect 1655 -1190 1705 -1160
rect 1915 -1175 1965 -1160
rect 1870 -1185 1965 -1175
rect 1450 -1225 1490 -1215
rect 1450 -1245 1460 -1225
rect 1480 -1230 1490 -1225
rect 1670 -1230 1685 -1190
rect 1870 -1205 1880 -1185
rect 1900 -1190 1965 -1185
rect 1900 -1205 1910 -1190
rect 1870 -1215 1910 -1205
rect 2015 -1200 2065 -1160
rect 2115 -1175 2165 -1160
rect 2215 -1175 2265 -1160
rect 2315 -1200 2365 -1160
rect 2415 -1175 2465 -1160
rect 2415 -1185 2510 -1175
rect 2415 -1190 2480 -1185
rect 2015 -1215 2365 -1200
rect 2470 -1205 2480 -1190
rect 2500 -1205 2510 -1185
rect 2470 -1215 2510 -1205
rect 1480 -1245 1685 -1230
rect 1450 -1255 1490 -1245
<< polycont >>
rect 2180 1460 2200 1480
rect 1540 1390 1560 1410
rect 1880 1415 1900 1435
rect 2480 1415 2500 1435
rect 1560 130 1580 150
rect 2180 145 2200 165
rect 1500 65 1520 85
rect 1460 -1180 1480 -1160
rect 1460 -1245 1480 -1225
rect 1880 -1205 1900 -1185
rect 2480 -1205 2500 -1185
<< locali >>
rect 2170 1485 2210 1490
rect 1435 1480 2210 1485
rect 1435 1465 2180 1480
rect 2170 1460 2180 1465
rect 2200 1460 2210 1480
rect 2170 1450 2210 1460
rect 1870 1435 1910 1445
rect 1435 1410 1570 1420
rect 1435 1400 1540 1410
rect 1530 1390 1540 1400
rect 1560 1390 1570 1410
rect 1530 1380 1570 1390
rect 1870 1415 1880 1435
rect 1900 1415 1910 1435
rect 1870 1385 1910 1415
rect 2470 1435 2510 1445
rect 2470 1415 2480 1435
rect 2500 1415 2510 1435
rect 2470 1385 2510 1415
rect 1590 1375 1630 1385
rect 1590 205 1600 1375
rect 1620 205 1630 1375
rect 1590 195 1630 205
rect 1690 1375 1780 1385
rect 1690 205 1700 1375
rect 1720 205 1750 1375
rect 1770 205 1780 1375
rect 1690 195 1780 205
rect 1820 1375 1910 1385
rect 1820 205 1830 1375
rect 1850 205 1880 1375
rect 1900 205 1910 1375
rect 1820 195 1910 205
rect 1970 1375 2010 1385
rect 1970 205 1980 1375
rect 2000 205 2010 1375
rect 1970 195 2010 205
rect 2070 1375 2110 1385
rect 2070 205 2080 1375
rect 2100 205 2110 1375
rect 2070 195 2110 205
rect 2170 1375 2210 1385
rect 2170 205 2180 1375
rect 2200 205 2210 1375
rect 2170 195 2210 205
rect 2270 1370 2310 1380
rect 2270 210 2280 1370
rect 2300 210 2310 1370
rect 2270 200 2310 210
rect 2370 1375 2410 1385
rect 2370 205 2380 1375
rect 2400 205 2410 1375
rect 2370 195 2410 205
rect 2470 1375 2560 1385
rect 2470 205 2480 1375
rect 2500 205 2530 1375
rect 2550 205 2560 1375
rect 2470 195 2560 205
rect 1550 150 1590 160
rect 1550 140 1560 150
rect 1435 130 1560 140
rect 1580 130 1590 150
rect 1435 120 1590 130
rect 1435 85 1530 95
rect 1435 75 1500 85
rect 1490 65 1500 75
rect 1520 65 1530 85
rect 1490 55 1530 65
rect 1610 35 1630 195
rect 1980 155 2000 195
rect 2170 165 2210 175
rect 2170 155 2180 165
rect 1980 145 2180 155
rect 2200 145 2210 165
rect 1980 135 2210 145
rect 1980 35 2000 135
rect 2380 105 2400 195
rect 2380 85 2585 105
rect 2380 35 2400 85
rect 1510 25 1550 35
rect 1510 -1145 1520 25
rect 1540 -1145 1550 25
rect 1435 -1160 1490 -1150
rect 1510 -1155 1550 -1145
rect 1610 25 1650 35
rect 1610 -1145 1620 25
rect 1640 -1145 1650 25
rect 1610 -1155 1650 -1145
rect 1710 25 1750 35
rect 1710 -1145 1720 25
rect 1740 -1145 1750 25
rect 1710 -1155 1750 -1145
rect 1820 25 1910 35
rect 1820 -1145 1830 25
rect 1850 -1145 1880 25
rect 1900 -1145 1910 25
rect 1820 -1155 1910 -1145
rect 1970 25 2010 35
rect 1970 -1145 1980 25
rect 2000 -1145 2010 25
rect 1970 -1155 2010 -1145
rect 2070 25 2110 35
rect 2070 -1145 2080 25
rect 2100 -1145 2110 25
rect 2070 -1155 2110 -1145
rect 2170 25 2210 35
rect 2170 -1145 2180 25
rect 2200 -1145 2210 25
rect 2170 -1155 2210 -1145
rect 2270 25 2310 35
rect 2270 -1145 2280 25
rect 2300 -1145 2310 25
rect 2270 -1155 2310 -1145
rect 2370 25 2410 35
rect 2370 -1145 2380 25
rect 2400 -1145 2410 25
rect 2370 -1155 2410 -1145
rect 2470 25 2560 35
rect 2470 -1145 2480 25
rect 2500 -1145 2530 25
rect 2550 -1145 2560 25
rect 2470 -1155 2560 -1145
rect 1435 -1170 1460 -1160
rect 1450 -1180 1460 -1170
rect 1480 -1180 1490 -1160
rect 1450 -1190 1490 -1180
rect 1435 -1225 1490 -1215
rect 1435 -1235 1460 -1225
rect 1450 -1245 1460 -1235
rect 1480 -1245 1490 -1225
rect 1450 -1255 1490 -1245
rect 1520 -1275 1540 -1155
rect 1720 -1235 1740 -1155
rect 1870 -1185 1910 -1155
rect 1870 -1205 1880 -1185
rect 1900 -1205 1910 -1185
rect 1870 -1215 1910 -1205
rect 2080 -1235 2100 -1155
rect 1720 -1255 2100 -1235
rect 2280 -1275 2300 -1155
rect 2470 -1185 2510 -1155
rect 2470 -1205 2480 -1185
rect 2500 -1205 2510 -1185
rect 2470 -1215 2510 -1205
rect 1520 -1295 2300 -1275
<< viali >>
rect 1700 205 1720 1375
rect 1750 205 1770 1375
rect 1830 205 1850 1375
rect 1880 205 1900 1375
rect 2180 205 2200 1375
rect 2480 205 2500 1375
rect 2530 205 2550 1375
rect 1830 -1145 1850 25
rect 1880 -1145 1900 25
rect 2180 -1145 2200 25
rect 2480 -1145 2500 25
rect 2530 -1145 2550 25
<< metal1 >>
rect 1435 1375 1785 1385
rect 1435 205 1700 1375
rect 1720 205 1750 1375
rect 1770 205 1785 1375
rect 1435 195 1785 205
rect 1815 1375 2585 1385
rect 1815 205 1830 1375
rect 1850 205 1880 1375
rect 1900 205 2180 1375
rect 2200 205 2480 1375
rect 2500 205 2530 1375
rect 2550 205 2585 1375
rect 1815 195 2585 205
rect 1435 25 2585 35
rect 1435 -1145 1830 25
rect 1850 -1145 1880 25
rect 1900 -1145 2180 25
rect 2200 -1145 2480 25
rect 2500 -1145 2530 25
rect 2550 -1145 2585 25
rect 1435 -1155 2585 -1145
<< labels >>
rlabel locali 2585 95 2585 95 3 Vout
rlabel locali 1435 130 1435 130 7 Vbn
rlabel locali 1435 -1225 1435 -1225 7 V1
rlabel locali 1435 -1160 1435 -1160 7 V2
rlabel locali 1435 85 1435 85 7 Vcn
rlabel locali 1435 1475 1435 1475 7 Vcp
rlabel locali 1435 1410 1435 1410 7 Vbp
rlabel metal1 1435 640 1435 640 7 VP
rlabel metal1 1435 -525 1435 -525 7 VN
<< end >>
