magic
tech sky130A
timestamp 1618804479
<< nwell >>
rect 1210 -150 3375 1090
rect 3135 -1625 3375 -150
<< nmos >>
rect 1330 -1605 1380 -405
rect 1430 -1605 1480 -405
rect 1530 -1605 1580 -405
rect 1630 -1605 1680 -405
rect 1730 -1605 1780 -405
rect 1830 -1605 1880 -405
rect 2110 -1605 2160 -405
rect 2210 -1605 2260 -405
rect 2310 -1605 2360 -405
rect 2410 -1605 2460 -405
rect 2510 -1605 2560 -405
rect 2740 -1605 2790 -405
rect 2970 -1605 3020 -405
<< pmos >>
rect 1330 -130 1380 1070
rect 1430 -130 1480 1070
rect 1530 -130 1580 1070
rect 1630 -130 1680 1070
rect 1730 -130 1780 1070
rect 1830 -130 1880 1070
rect 1930 -130 1980 1070
rect 2210 -130 2260 1070
rect 2310 -130 2360 1070
rect 2410 -130 2460 1070
rect 2510 -130 2560 1070
rect 2610 -130 2660 1070
rect 2710 -130 2760 1070
rect 2810 -130 2860 1070
rect 3040 -130 3090 1070
rect 3140 -130 3190 1070
rect 3255 -1605 3305 -405
<< ndiff >>
rect 1280 -420 1330 -405
rect 1280 -1590 1295 -420
rect 1315 -1590 1330 -420
rect 1280 -1605 1330 -1590
rect 1380 -420 1430 -405
rect 1380 -1590 1395 -420
rect 1415 -1590 1430 -420
rect 1380 -1605 1430 -1590
rect 1480 -420 1530 -405
rect 1480 -1590 1495 -420
rect 1515 -1590 1530 -420
rect 1480 -1605 1530 -1590
rect 1580 -420 1630 -405
rect 1580 -1590 1595 -420
rect 1615 -1590 1630 -420
rect 1580 -1605 1630 -1590
rect 1680 -420 1730 -405
rect 1680 -1590 1695 -420
rect 1715 -1590 1730 -420
rect 1680 -1605 1730 -1590
rect 1780 -420 1830 -405
rect 1780 -1590 1795 -420
rect 1815 -1590 1830 -420
rect 1780 -1605 1830 -1590
rect 1880 -420 1930 -405
rect 1880 -1590 1895 -420
rect 1915 -1590 1930 -420
rect 1880 -1605 1930 -1590
rect 2060 -420 2110 -405
rect 2060 -1590 2075 -420
rect 2095 -1590 2110 -420
rect 2060 -1605 2110 -1590
rect 2160 -420 2210 -405
rect 2160 -1590 2175 -420
rect 2195 -1590 2210 -420
rect 2160 -1605 2210 -1590
rect 2260 -420 2310 -405
rect 2260 -1590 2275 -420
rect 2295 -1590 2310 -420
rect 2260 -1605 2310 -1590
rect 2360 -420 2410 -405
rect 2360 -1590 2375 -420
rect 2395 -1590 2410 -420
rect 2360 -1605 2410 -1590
rect 2460 -420 2510 -405
rect 2460 -1590 2475 -420
rect 2495 -1590 2510 -420
rect 2460 -1605 2510 -1590
rect 2560 -420 2610 -405
rect 2560 -1590 2575 -420
rect 2595 -1590 2610 -420
rect 2560 -1605 2610 -1590
rect 2690 -420 2740 -405
rect 2690 -1590 2705 -420
rect 2725 -1590 2740 -420
rect 2690 -1605 2740 -1590
rect 2790 -420 2840 -405
rect 2790 -1590 2805 -420
rect 2825 -1590 2840 -420
rect 2790 -1605 2840 -1590
rect 2920 -420 2970 -405
rect 2920 -1590 2935 -420
rect 2955 -1590 2970 -420
rect 2920 -1605 2970 -1590
rect 3020 -420 3070 -405
rect 3020 -1590 3035 -420
rect 3055 -1590 3070 -420
rect 3020 -1605 3070 -1590
<< pdiff >>
rect 1280 1055 1330 1070
rect 1280 -115 1295 1055
rect 1315 -115 1330 1055
rect 1280 -130 1330 -115
rect 1380 1055 1430 1070
rect 1380 -115 1395 1055
rect 1415 -115 1430 1055
rect 1380 -130 1430 -115
rect 1480 1055 1530 1070
rect 1480 -115 1495 1055
rect 1515 -115 1530 1055
rect 1480 -130 1530 -115
rect 1580 1055 1630 1070
rect 1580 -115 1595 1055
rect 1615 -115 1630 1055
rect 1580 -130 1630 -115
rect 1680 1055 1730 1070
rect 1680 -115 1695 1055
rect 1715 -115 1730 1055
rect 1680 -130 1730 -115
rect 1780 1055 1830 1070
rect 1780 -115 1795 1055
rect 1815 -115 1830 1055
rect 1780 -130 1830 -115
rect 1880 1055 1930 1070
rect 1880 -115 1895 1055
rect 1915 -115 1930 1055
rect 1880 -130 1930 -115
rect 1980 1055 2030 1070
rect 1980 -115 1995 1055
rect 2015 -115 2030 1055
rect 1980 -130 2030 -115
rect 2160 1055 2210 1070
rect 2160 -115 2175 1055
rect 2195 -115 2210 1055
rect 2160 -130 2210 -115
rect 2260 1055 2310 1070
rect 2260 -115 2275 1055
rect 2295 -115 2310 1055
rect 2260 -130 2310 -115
rect 2360 1055 2410 1070
rect 2360 -115 2375 1055
rect 2395 -115 2410 1055
rect 2360 -130 2410 -115
rect 2460 1055 2510 1070
rect 2460 -115 2475 1055
rect 2495 -115 2510 1055
rect 2460 -130 2510 -115
rect 2560 1055 2610 1070
rect 2560 -115 2575 1055
rect 2595 -115 2610 1055
rect 2560 -130 2610 -115
rect 2660 1055 2710 1070
rect 2660 -115 2675 1055
rect 2695 -115 2710 1055
rect 2660 -130 2710 -115
rect 2760 1055 2810 1070
rect 2760 -115 2775 1055
rect 2795 -115 2810 1055
rect 2760 -130 2810 -115
rect 2860 1055 2910 1070
rect 2860 -115 2875 1055
rect 2895 -115 2910 1055
rect 2860 -130 2910 -115
rect 2990 1055 3040 1070
rect 2990 -115 3005 1055
rect 3025 -115 3040 1055
rect 2990 -130 3040 -115
rect 3090 1055 3140 1070
rect 3090 -115 3105 1055
rect 3125 -115 3140 1055
rect 3090 -130 3140 -115
rect 3190 1055 3240 1070
rect 3190 -115 3205 1055
rect 3225 -115 3240 1055
rect 3190 -130 3240 -115
rect 3205 -420 3255 -405
rect 3205 -1590 3220 -420
rect 3240 -1590 3255 -420
rect 3205 -1605 3255 -1590
rect 3305 -420 3355 -405
rect 3305 -1590 3320 -420
rect 3340 -1590 3355 -420
rect 3305 -1605 3355 -1590
<< ndiffc >>
rect 1295 -1590 1315 -420
rect 1395 -1590 1415 -420
rect 1495 -1590 1515 -420
rect 1595 -1590 1615 -420
rect 1695 -1590 1715 -420
rect 1795 -1590 1815 -420
rect 1895 -1590 1915 -420
rect 2075 -1590 2095 -420
rect 2175 -1590 2195 -420
rect 2275 -1590 2295 -420
rect 2375 -1590 2395 -420
rect 2475 -1590 2495 -420
rect 2575 -1590 2595 -420
rect 2705 -1590 2725 -420
rect 2805 -1590 2825 -420
rect 2935 -1590 2955 -420
rect 3035 -1590 3055 -420
<< pdiffc >>
rect 1295 -115 1315 1055
rect 1395 -115 1415 1055
rect 1495 -115 1515 1055
rect 1595 -115 1615 1055
rect 1695 -115 1715 1055
rect 1795 -115 1815 1055
rect 1895 -115 1915 1055
rect 1995 -115 2015 1055
rect 2175 -115 2195 1055
rect 2275 -115 2295 1055
rect 2375 -115 2395 1055
rect 2475 -115 2495 1055
rect 2575 -115 2595 1055
rect 2675 -115 2695 1055
rect 2775 -115 2795 1055
rect 2875 -115 2895 1055
rect 3005 -115 3025 1055
rect 3105 -115 3125 1055
rect 3205 -115 3225 1055
rect 3220 -1590 3240 -420
rect 3320 -1590 3340 -420
<< psubdiff >>
rect 1230 -420 1280 -405
rect 1230 -1590 1245 -420
rect 1265 -1590 1280 -420
rect 1230 -1605 1280 -1590
rect 1930 -420 1980 -405
rect 1930 -1590 1945 -420
rect 1965 -1590 1980 -420
rect 1930 -1605 1980 -1590
rect 2010 -420 2060 -405
rect 2010 -1590 2025 -420
rect 2045 -1590 2060 -420
rect 2010 -1605 2060 -1590
rect 2610 -420 2660 -405
rect 2610 -1590 2625 -420
rect 2645 -1590 2660 -420
rect 2610 -1605 2660 -1590
rect 2840 -420 2890 -405
rect 2840 -1590 2855 -420
rect 2875 -1590 2890 -420
rect 2840 -1605 2890 -1590
rect 3070 -420 3120 -405
rect 3070 -1590 3085 -420
rect 3105 -1590 3120 -420
rect 3070 -1605 3120 -1590
<< nsubdiff >>
rect 1230 1055 1280 1070
rect 1230 -115 1245 1055
rect 1265 -115 1280 1055
rect 1230 -130 1280 -115
rect 2030 1055 2080 1070
rect 2030 -115 2045 1055
rect 2065 -115 2080 1055
rect 2030 -130 2080 -115
rect 2110 1055 2160 1070
rect 2110 -115 2125 1055
rect 2145 -115 2160 1055
rect 2110 -130 2160 -115
rect 2910 1055 2960 1070
rect 2910 -115 2925 1055
rect 2945 -115 2960 1055
rect 2910 -130 2960 -115
rect 3240 1055 3290 1070
rect 3240 -115 3255 1055
rect 3275 -115 3290 1055
rect 3240 -130 3290 -115
rect 3155 -420 3205 -405
rect 3155 -1590 3170 -420
rect 3190 -1590 3205 -420
rect 3155 -1605 3205 -1590
<< psubdiffcont >>
rect 1245 -1590 1265 -420
rect 1945 -1590 1965 -420
rect 2025 -1590 2045 -420
rect 2625 -1590 2645 -420
rect 2855 -1590 2875 -420
rect 3085 -1590 3105 -420
<< nsubdiffcont >>
rect 1245 -115 1265 1055
rect 2045 -115 2065 1055
rect 2125 -115 2145 1055
rect 2925 -115 2945 1055
rect 3255 -115 3275 1055
rect 3170 -1590 3190 -420
<< poly >>
rect 1285 1115 1325 1125
rect 1285 1095 1295 1115
rect 1315 1100 1325 1115
rect 1830 1110 2360 1125
rect 1830 1100 1880 1110
rect 1315 1095 1380 1100
rect 1285 1085 1380 1095
rect 1330 1070 1380 1085
rect 1430 1085 1880 1100
rect 2310 1100 2360 1110
rect 2860 1115 2900 1125
rect 2860 1100 2870 1115
rect 2310 1085 2760 1100
rect 1430 1070 1480 1085
rect 1530 1070 1580 1085
rect 1630 1070 1680 1085
rect 1730 1070 1780 1085
rect 1830 1070 1880 1085
rect 1930 1070 1980 1085
rect 2210 1070 2260 1085
rect 2310 1070 2360 1085
rect 2410 1070 2460 1085
rect 2510 1070 2560 1085
rect 2610 1070 2660 1085
rect 2710 1070 2760 1085
rect 2810 1095 2870 1100
rect 2890 1095 2900 1115
rect 2810 1085 2900 1095
rect 3000 1115 3040 1125
rect 3000 1095 3010 1115
rect 3030 1100 3040 1115
rect 3030 1095 3190 1100
rect 3000 1085 3190 1095
rect 2810 1070 2860 1085
rect 3040 1070 3090 1085
rect 3140 1070 3190 1085
rect 1330 -145 1380 -130
rect 1430 -145 1480 -130
rect 1530 -145 1580 -130
rect 1630 -145 1680 -130
rect 1730 -145 1780 -130
rect 1830 -145 1880 -130
rect 1930 -145 1980 -130
rect 2210 -145 2260 -130
rect 2310 -145 2360 -130
rect 2410 -145 2460 -130
rect 2510 -145 2560 -130
rect 2610 -145 2660 -130
rect 2710 -145 2760 -130
rect 2810 -145 2860 -130
rect 3040 -145 3090 -130
rect 3140 -145 3190 -130
rect 1635 -155 1675 -145
rect 1635 -175 1645 -155
rect 1665 -175 1675 -155
rect 1930 -155 2020 -145
rect 1930 -160 1990 -155
rect 1635 -185 1675 -175
rect 1980 -175 1990 -160
rect 2010 -175 2020 -155
rect 1980 -185 2020 -175
rect 2170 -155 2260 -145
rect 2170 -175 2180 -155
rect 2200 -160 2260 -155
rect 2200 -175 2210 -160
rect 2170 -185 2210 -175
rect 3205 -170 3245 -160
rect 3205 -185 3215 -170
rect 1660 -210 1675 -185
rect 2880 -190 3215 -185
rect 3235 -190 3245 -170
rect 2880 -200 3245 -190
rect 2880 -210 2895 -200
rect 1660 -225 2895 -210
rect 2980 -240 3245 -230
rect 2980 -245 3215 -240
rect 2980 -250 2995 -245
rect 2235 -265 2995 -250
rect 3205 -260 3215 -245
rect 3235 -260 3245 -240
rect 2235 -350 2250 -265
rect 3205 -270 3245 -260
rect 3205 -310 3245 -300
rect 2720 -325 3215 -310
rect 2415 -350 2455 -340
rect 2720 -350 2735 -325
rect 3205 -330 3215 -325
rect 3235 -330 3245 -310
rect 3205 -340 3245 -330
rect 1290 -360 1330 -350
rect 1290 -380 1300 -360
rect 1320 -375 1330 -360
rect 1880 -360 1920 -350
rect 1880 -375 1890 -360
rect 1320 -380 1380 -375
rect 1290 -390 1380 -380
rect 1830 -380 1890 -375
rect 1910 -380 1920 -360
rect 1830 -390 1920 -380
rect 2070 -360 2110 -350
rect 2070 -380 2080 -360
rect 2100 -375 2110 -360
rect 2215 -360 2255 -350
rect 2100 -380 2160 -375
rect 2070 -390 2160 -380
rect 2215 -380 2225 -360
rect 2245 -380 2255 -360
rect 2415 -370 2425 -350
rect 2445 -370 2455 -350
rect 2415 -380 2455 -370
rect 2560 -360 2600 -350
rect 2560 -375 2570 -360
rect 2510 -380 2570 -375
rect 2590 -380 2600 -360
rect 2215 -390 2255 -380
rect 1330 -405 1380 -390
rect 1430 -405 1480 -390
rect 1530 -405 1580 -390
rect 1630 -405 1680 -390
rect 1730 -405 1780 -390
rect 1830 -405 1880 -390
rect 2110 -405 2160 -390
rect 2210 -405 2260 -390
rect 2310 -395 2460 -380
rect 2310 -405 2360 -395
rect 2410 -405 2460 -395
rect 2510 -390 2600 -380
rect 2700 -360 2740 -350
rect 2700 -380 2710 -360
rect 2730 -375 2740 -360
rect 3305 -360 3345 -350
rect 3305 -375 3315 -360
rect 2730 -380 2790 -375
rect 2700 -390 2790 -380
rect 3255 -380 3315 -375
rect 3335 -380 3345 -360
rect 3255 -390 3345 -380
rect 2510 -405 2560 -390
rect 2740 -405 2790 -390
rect 2970 -405 3020 -390
rect 3255 -405 3305 -390
rect 1330 -1620 1380 -1605
rect 1430 -1645 1480 -1605
rect 1530 -1645 1580 -1605
rect 1630 -1645 1680 -1605
rect 1730 -1645 1780 -1605
rect 1830 -1620 1880 -1605
rect 2110 -1620 2160 -1605
rect 2210 -1645 2260 -1605
rect 2310 -1620 2360 -1605
rect 2410 -1620 2460 -1605
rect 2510 -1620 2560 -1605
rect 2740 -1620 2790 -1605
rect 2970 -1645 3020 -1605
rect 3255 -1620 3305 -1605
rect 1430 -1660 3020 -1645
<< polycont >>
rect 1295 1095 1315 1115
rect 2870 1095 2890 1115
rect 3010 1095 3030 1115
rect 1645 -175 1665 -155
rect 1990 -175 2010 -155
rect 2180 -175 2200 -155
rect 3215 -190 3235 -170
rect 3215 -260 3235 -240
rect 3215 -330 3235 -310
rect 1300 -380 1320 -360
rect 1890 -380 1910 -360
rect 2080 -380 2100 -360
rect 2225 -380 2245 -360
rect 2425 -370 2445 -350
rect 2570 -380 2590 -360
rect 2710 -380 2730 -360
rect 3315 -380 3335 -360
<< locali >>
rect 1285 1115 1325 1125
rect 1285 1095 1295 1115
rect 1315 1095 1325 1115
rect 1285 1065 1325 1095
rect 1395 1100 1815 1120
rect 1395 1065 1415 1100
rect 1595 1065 1615 1100
rect 1795 1065 1815 1100
rect 2385 1100 2795 1120
rect 2385 1065 2405 1100
rect 2575 1065 2595 1100
rect 2775 1065 2795 1100
rect 2860 1115 2900 1125
rect 2860 1095 2870 1115
rect 2890 1095 2900 1115
rect 2860 1085 2900 1095
rect 2865 1065 2900 1085
rect 3000 1115 3040 1125
rect 3000 1095 3010 1115
rect 3030 1095 3040 1115
rect 3000 1085 3040 1095
rect 3000 1065 3035 1085
rect 1235 1055 1325 1065
rect 1235 -115 1245 1055
rect 1265 -115 1295 1055
rect 1315 -115 1325 1055
rect 1235 -125 1325 -115
rect 1385 1055 1425 1065
rect 1385 -115 1395 1055
rect 1415 -115 1425 1055
rect 1385 -125 1425 -115
rect 1485 1055 1525 1065
rect 1485 -115 1495 1055
rect 1515 -115 1525 1055
rect 1485 -125 1525 -115
rect 1585 1055 1625 1065
rect 1585 -115 1595 1055
rect 1615 -115 1625 1055
rect 1585 -125 1625 -115
rect 1685 1055 1725 1065
rect 1685 -115 1695 1055
rect 1715 -115 1725 1055
rect 1685 -125 1725 -115
rect 1785 1055 1825 1065
rect 1785 -115 1795 1055
rect 1815 -115 1825 1055
rect 1785 -125 1825 -115
rect 1885 1055 1925 1065
rect 1885 -115 1895 1055
rect 1915 -115 1925 1055
rect 1885 -125 1925 -115
rect 1495 -145 1515 -125
rect 1695 -145 1715 -125
rect 1210 -155 1715 -145
rect 1210 -165 1645 -155
rect 1635 -175 1645 -165
rect 1665 -165 1715 -155
rect 1665 -175 1675 -165
rect 1635 -185 1675 -175
rect 1905 -285 1925 -125
rect 1985 1055 2075 1065
rect 1985 -115 1995 1055
rect 2015 -115 2045 1055
rect 2065 -115 2075 1055
rect 1985 -125 2075 -115
rect 2115 1055 2205 1065
rect 2115 -115 2125 1055
rect 2145 -115 2175 1055
rect 2195 -115 2205 1055
rect 2115 -125 2205 -115
rect 2265 1055 2305 1065
rect 2265 -115 2275 1055
rect 2295 -115 2305 1055
rect 2265 -125 2305 -115
rect 2365 1055 2405 1065
rect 2365 -115 2375 1055
rect 2395 -115 2405 1055
rect 2365 -125 2405 -115
rect 2465 1055 2505 1065
rect 2465 -115 2475 1055
rect 2495 -115 2505 1055
rect 2465 -125 2505 -115
rect 2565 1055 2605 1065
rect 2565 -115 2575 1055
rect 2595 -115 2605 1055
rect 2565 -125 2605 -115
rect 2665 1055 2705 1065
rect 2665 -115 2675 1055
rect 2695 -115 2705 1055
rect 2665 -125 2705 -115
rect 2765 1055 2805 1065
rect 2765 -115 2775 1055
rect 2795 -115 2805 1055
rect 2765 -125 2805 -115
rect 2865 1055 2955 1065
rect 2865 -115 2875 1055
rect 2895 -115 2925 1055
rect 2945 -115 2955 1055
rect 2865 -125 2955 -115
rect 2995 1055 3035 1065
rect 2995 -115 3005 1055
rect 3025 -115 3035 1055
rect 2995 -125 3035 -115
rect 3095 1055 3135 1065
rect 3095 -115 3105 1055
rect 3125 -115 3135 1055
rect 3095 -125 3135 -115
rect 3195 1055 3285 1065
rect 3195 -115 3205 1055
rect 3225 -115 3255 1055
rect 3275 -115 3285 1055
rect 3195 -125 3285 -115
rect 1985 -145 2020 -125
rect 1980 -155 2020 -145
rect 1980 -175 1990 -155
rect 2010 -175 2020 -155
rect 1980 -185 2020 -175
rect 2170 -145 2205 -125
rect 2170 -155 2210 -145
rect 2170 -175 2180 -155
rect 2200 -175 2210 -155
rect 2170 -185 2210 -175
rect 2285 -190 2305 -125
rect 2475 -145 2495 -125
rect 2675 -145 2695 -125
rect 2475 -165 2720 -145
rect 3005 -150 3025 -125
rect 2285 -210 2485 -190
rect 1905 -305 2235 -285
rect 2215 -350 2235 -305
rect 2465 -340 2485 -210
rect 2415 -350 2485 -340
rect 2700 -350 2720 -165
rect 2945 -170 3025 -150
rect 3105 -145 3125 -125
rect 3105 -165 3180 -145
rect 1290 -360 1330 -350
rect 1290 -380 1300 -360
rect 1320 -380 1330 -360
rect 1880 -360 1920 -350
rect 1290 -390 1330 -380
rect 1395 -390 1815 -370
rect 1880 -380 1890 -360
rect 1910 -380 1920 -360
rect 1880 -390 1920 -380
rect 1290 -410 1325 -390
rect 1395 -410 1415 -390
rect 1595 -410 1615 -390
rect 1795 -410 1815 -390
rect 1885 -410 1920 -390
rect 2070 -360 2110 -350
rect 2070 -380 2080 -360
rect 2100 -380 2110 -360
rect 2215 -360 2255 -350
rect 2215 -370 2225 -360
rect 2070 -390 2110 -380
rect 2185 -380 2225 -370
rect 2245 -380 2255 -360
rect 2415 -370 2425 -350
rect 2445 -370 2485 -350
rect 2415 -380 2485 -370
rect 2185 -390 2255 -380
rect 2070 -410 2105 -390
rect 2185 -410 2205 -390
rect 2465 -410 2485 -380
rect 2560 -360 2600 -350
rect 2560 -380 2570 -360
rect 2590 -380 2600 -360
rect 2560 -390 2600 -380
rect 2565 -410 2600 -390
rect 2700 -360 2740 -350
rect 2700 -380 2710 -360
rect 2730 -380 2740 -360
rect 2700 -390 2740 -380
rect 2700 -410 2735 -390
rect 2945 -410 2965 -170
rect 3160 -410 3180 -165
rect 3205 -170 3375 -160
rect 3205 -190 3215 -170
rect 3235 -180 3375 -170
rect 3235 -190 3245 -180
rect 3205 -200 3245 -190
rect 3205 -240 3375 -230
rect 3205 -260 3215 -240
rect 3235 -250 3375 -240
rect 3235 -260 3245 -250
rect 3205 -270 3245 -260
rect 3205 -310 3375 -300
rect 3205 -330 3215 -310
rect 3235 -320 3375 -310
rect 3235 -330 3245 -320
rect 3205 -340 3245 -330
rect 3305 -360 3345 -350
rect 3305 -380 3315 -360
rect 3335 -370 3345 -360
rect 3335 -380 3375 -370
rect 3305 -390 3375 -380
rect 3310 -410 3345 -390
rect 1235 -420 1325 -410
rect 1235 -1590 1245 -420
rect 1265 -1590 1295 -420
rect 1315 -1590 1325 -420
rect 1235 -1600 1325 -1590
rect 1385 -420 1425 -410
rect 1385 -1590 1395 -420
rect 1415 -1590 1425 -420
rect 1385 -1600 1425 -1590
rect 1485 -420 1525 -410
rect 1485 -1590 1495 -420
rect 1515 -1590 1525 -420
rect 1485 -1600 1525 -1590
rect 1585 -420 1625 -410
rect 1585 -1590 1595 -420
rect 1615 -1590 1625 -420
rect 1585 -1600 1625 -1590
rect 1685 -420 1725 -410
rect 1685 -1590 1695 -420
rect 1715 -1590 1725 -420
rect 1685 -1600 1725 -1590
rect 1785 -420 1825 -410
rect 1785 -1590 1795 -420
rect 1815 -1590 1825 -420
rect 1785 -1600 1825 -1590
rect 1885 -420 1975 -410
rect 1885 -1590 1895 -420
rect 1915 -1590 1945 -420
rect 1965 -1590 1975 -420
rect 1885 -1600 1975 -1590
rect 2015 -420 2105 -410
rect 2015 -1590 2025 -420
rect 2045 -1590 2075 -420
rect 2095 -1590 2105 -420
rect 2015 -1600 2105 -1590
rect 2165 -420 2205 -410
rect 2165 -1590 2175 -420
rect 2195 -1590 2205 -420
rect 2165 -1600 2205 -1590
rect 2265 -420 2305 -410
rect 2265 -1590 2275 -420
rect 2295 -1590 2305 -420
rect 2265 -1600 2305 -1590
rect 2365 -420 2405 -410
rect 2365 -1590 2375 -420
rect 2395 -1590 2405 -420
rect 2365 -1600 2405 -1590
rect 2465 -420 2505 -410
rect 2465 -1590 2475 -420
rect 2495 -1590 2505 -420
rect 2465 -1600 2505 -1590
rect 2565 -420 2655 -410
rect 2565 -1590 2575 -420
rect 2595 -1590 2625 -420
rect 2645 -1590 2655 -420
rect 2565 -1600 2655 -1590
rect 2695 -420 2735 -410
rect 2695 -1590 2705 -420
rect 2725 -1590 2735 -420
rect 2695 -1600 2735 -1590
rect 2795 -420 2885 -410
rect 2795 -1590 2805 -420
rect 2825 -1590 2855 -420
rect 2875 -1590 2885 -420
rect 2795 -1600 2885 -1590
rect 2925 -420 2965 -410
rect 2925 -1590 2935 -420
rect 2955 -1590 2965 -420
rect 2925 -1600 2965 -1590
rect 3025 -420 3115 -410
rect 3025 -1590 3035 -420
rect 3055 -1590 3085 -420
rect 3105 -1590 3115 -420
rect 3025 -1600 3115 -1590
rect 3160 -420 3250 -410
rect 3160 -1590 3170 -420
rect 3190 -1590 3220 -420
rect 3240 -1590 3250 -420
rect 3160 -1600 3250 -1590
rect 3310 -420 3350 -410
rect 3310 -1590 3320 -420
rect 3340 -1590 3350 -420
rect 3310 -1600 3350 -1590
rect 1495 -1660 1515 -1600
rect 1695 -1660 1715 -1600
rect 2375 -1620 2395 -1600
rect 2795 -1620 2815 -1600
rect 2375 -1640 2815 -1620
rect 3310 -1660 3330 -1600
rect 1495 -1680 3330 -1660
<< viali >>
rect 1245 -115 1265 1055
rect 1295 -115 1315 1055
rect 1395 -115 1415 1055
rect 1595 -115 1615 1055
rect 1795 -115 1815 1055
rect 1995 -115 2015 1055
rect 2045 -115 2065 1055
rect 2125 -115 2145 1055
rect 2175 -115 2195 1055
rect 2375 -115 2395 1055
rect 2575 -115 2595 1055
rect 2775 -115 2795 1055
rect 2875 -115 2895 1055
rect 2925 -115 2945 1055
rect 3205 -115 3225 1055
rect 3255 -115 3275 1055
rect 1245 -1590 1265 -420
rect 1295 -1590 1315 -420
rect 1395 -1590 1415 -420
rect 1595 -1590 1615 -420
rect 1795 -1590 1815 -420
rect 1895 -1590 1915 -420
rect 1945 -1590 1965 -420
rect 2025 -1590 2045 -420
rect 2075 -1590 2095 -420
rect 2275 -1590 2295 -420
rect 2575 -1590 2595 -420
rect 2625 -1590 2645 -420
rect 3035 -1590 3055 -420
rect 3085 -1590 3105 -420
<< metal1 >>
rect 1210 1055 3375 1065
rect 1210 -115 1245 1055
rect 1265 -115 1295 1055
rect 1315 -115 1395 1055
rect 1415 -115 1595 1055
rect 1615 -115 1795 1055
rect 1815 -115 1995 1055
rect 2015 -115 2045 1055
rect 2065 -115 2125 1055
rect 2145 -115 2175 1055
rect 2195 -115 2375 1055
rect 2395 -115 2575 1055
rect 2595 -115 2775 1055
rect 2795 -115 2875 1055
rect 2895 -115 2925 1055
rect 2945 -115 3205 1055
rect 3225 -115 3255 1055
rect 3275 -115 3375 1055
rect 1210 -125 3375 -115
rect 1210 -420 3375 -410
rect 1210 -1590 1245 -420
rect 1265 -1590 1295 -420
rect 1315 -1590 1395 -420
rect 1415 -1590 1595 -420
rect 1615 -1590 1795 -420
rect 1815 -1590 1895 -420
rect 1915 -1590 1945 -420
rect 1965 -1590 2025 -420
rect 2045 -1590 2075 -420
rect 2095 -1590 2275 -420
rect 2295 -1590 2575 -420
rect 2595 -1590 2625 -420
rect 2645 -1590 3035 -420
rect 3055 -1590 3085 -420
rect 3105 -1590 3375 -420
rect 1210 -1600 3375 -1590
<< labels >>
rlabel locali 1210 -155 1210 -155 7 Vb
rlabel locali 3375 -240 3375 -240 3 Vbn
rlabel locali 3375 -310 3375 -310 3 Vcn
rlabel metal1 1210 -945 1210 -945 7 VN
rlabel metal1 1210 370 1210 370 7 VP
rlabel locali 3375 -380 3375 -380 3 Vcp
<< end >>
