magic
tech sky130A
timestamp 1616037287
<< error_p >>
rect 1044 603 1050 606
rect 1264 603 1270 606
rect 1484 603 1490 606
rect 1027 600 1053 603
rect 1247 600 1273 603
rect 1467 600 1493 603
rect 1024 597 1056 600
rect 1024 594 1033 597
rect 1030 523 1033 594
rect 1047 594 1056 597
rect 1244 597 1276 600
rect 1244 594 1253 597
rect 1047 523 1053 594
rect 1030 520 1053 523
rect 1250 523 1253 594
rect 1267 594 1276 597
rect 1464 597 1496 600
rect 1464 594 1473 597
rect 1267 523 1273 594
rect 1250 520 1273 523
rect 1470 523 1473 594
rect 1487 594 1496 597
rect 1487 523 1493 594
rect 1470 520 1493 523
rect 1044 517 1053 520
rect 1264 517 1273 520
rect 1484 517 1493 520
rect 1044 514 1050 517
rect 1264 514 1270 517
rect 1484 514 1490 517
<< nwell >>
rect 690 460 1660 660
<< nmos >>
rect 850 200 900 320
<< pmos >>
rect 850 500 900 620
rect 960 500 1010 620
rect 1070 500 1120 620
rect 1180 500 1230 620
rect 1290 500 1340 620
rect 1400 500 1450 620
rect 1510 500 1560 620
<< ndiff >>
rect 790 300 850 320
rect 790 220 810 300
rect 830 220 850 300
rect 790 200 850 220
rect 900 300 960 320
rect 900 220 920 300
rect 940 220 960 300
rect 900 200 960 220
<< pdiff >>
rect 790 600 850 620
rect 790 520 810 600
rect 830 520 850 600
rect 790 500 850 520
rect 900 600 960 620
rect 900 520 920 600
rect 940 520 960 600
rect 900 500 960 520
rect 1010 600 1070 620
rect 1010 520 1030 600
rect 1050 520 1070 600
rect 1010 500 1070 520
rect 1120 600 1180 620
rect 1120 520 1140 600
rect 1160 520 1180 600
rect 1120 500 1180 520
rect 1230 600 1290 620
rect 1230 520 1250 600
rect 1270 520 1290 600
rect 1230 500 1290 520
rect 1340 600 1400 620
rect 1340 520 1360 600
rect 1380 520 1400 600
rect 1340 500 1400 520
rect 1450 600 1510 620
rect 1450 520 1470 600
rect 1490 520 1510 600
rect 1450 500 1510 520
rect 1560 600 1620 620
rect 1560 520 1580 600
rect 1600 520 1620 600
rect 1560 500 1620 520
<< ndiffc >>
rect 810 220 830 300
rect 920 220 940 300
<< pdiffc >>
rect 810 520 830 600
rect 920 520 940 600
rect 1030 520 1050 600
rect 1140 520 1160 600
rect 1250 520 1270 600
rect 1360 520 1380 600
rect 1470 520 1490 600
rect 1580 520 1600 600
<< psubdiff >>
rect 730 300 790 320
rect 730 220 750 300
rect 770 220 790 300
rect 730 200 790 220
<< nsubdiff >>
rect 730 600 790 620
rect 730 520 750 600
rect 770 520 790 600
rect 730 500 790 520
<< psubdiffcont >>
rect 750 220 770 300
<< nsubdiffcont >>
rect 750 520 770 600
<< poly >>
rect 850 700 910 710
rect 850 660 860 700
rect 900 660 910 700
rect 850 650 910 660
rect 960 700 1020 710
rect 960 660 970 700
rect 1010 660 1020 700
rect 960 650 1020 660
rect 1070 700 1130 710
rect 1070 660 1080 700
rect 1120 660 1130 700
rect 1070 650 1130 660
rect 1180 700 1240 710
rect 1180 660 1190 700
rect 1230 660 1240 700
rect 1180 650 1240 660
rect 1290 700 1350 710
rect 1290 660 1300 700
rect 1340 660 1350 700
rect 1290 650 1350 660
rect 1400 700 1460 710
rect 1400 660 1410 700
rect 1450 660 1460 700
rect 1400 650 1460 660
rect 1510 700 1570 710
rect 1510 660 1520 700
rect 1560 660 1570 700
rect 1510 650 1570 660
rect 850 620 900 650
rect 960 620 1010 650
rect 1070 620 1120 650
rect 1180 620 1230 650
rect 1290 620 1340 650
rect 1400 620 1450 650
rect 1510 620 1560 650
rect 850 470 900 500
rect 960 470 1010 500
rect 1070 470 1120 500
rect 1180 470 1230 500
rect 1290 470 1340 500
rect 1400 470 1450 500
rect 1510 470 1560 500
rect 850 320 900 350
rect 850 170 900 200
<< polycont >>
rect 860 660 900 700
rect 970 660 1010 700
rect 1080 660 1120 700
rect 1190 660 1230 700
rect 1300 660 1340 700
rect 1410 660 1450 700
rect 1520 660 1560 700
<< locali >>
rect 850 700 1570 710
rect 850 660 860 700
rect 900 670 970 700
rect 900 660 910 670
rect 850 650 910 660
rect 960 660 970 670
rect 1010 670 1080 700
rect 1010 660 1020 670
rect 960 650 1020 660
rect 1070 660 1080 670
rect 1120 670 1190 700
rect 1120 660 1130 670
rect 1070 650 1130 660
rect 1180 660 1190 670
rect 1230 670 1300 700
rect 1230 660 1240 670
rect 1180 650 1240 660
rect 1290 660 1300 670
rect 1340 670 1410 700
rect 1340 660 1350 670
rect 1290 650 1350 660
rect 1400 660 1410 670
rect 1450 670 1520 700
rect 1450 660 1460 670
rect 1400 650 1460 660
rect 1510 660 1520 670
rect 1560 660 1570 700
rect 1510 650 1570 660
rect 740 600 840 610
rect 740 520 750 600
rect 770 520 810 600
rect 830 520 840 600
rect 740 510 840 520
rect 910 600 950 610
rect 910 520 920 600
rect 940 520 950 600
rect 910 510 950 520
rect 1020 600 1060 610
rect 1020 520 1030 600
rect 1050 520 1060 600
rect 1020 510 1060 520
rect 1130 600 1170 610
rect 1130 520 1140 600
rect 1160 520 1170 600
rect 1130 510 1170 520
rect 1240 600 1280 610
rect 1240 520 1250 600
rect 1270 520 1280 600
rect 1240 510 1280 520
rect 1350 600 1390 610
rect 1350 520 1360 600
rect 1380 520 1390 600
rect 1350 510 1390 520
rect 1460 600 1500 610
rect 1460 520 1470 600
rect 1490 520 1500 600
rect 1460 510 1500 520
rect 1570 600 1610 610
rect 1570 520 1580 600
rect 1600 520 1610 600
rect 1570 510 1610 520
rect 920 450 940 510
rect 1140 450 1160 510
rect 1360 450 1380 510
rect 1580 450 1600 510
rect 920 430 1600 450
rect 740 300 840 310
rect 740 220 750 300
rect 770 220 810 300
rect 830 220 840 300
rect 740 210 840 220
rect 910 300 950 310
rect 910 220 920 300
rect 940 220 950 300
rect 910 210 950 220
<< viali >>
rect 1030 520 1050 600
rect 1250 520 1270 600
rect 1470 520 1490 600
<< end >>
