* SPICE3 file created from AND.ext - technology: sky130A

.subckt inverter VP VN A Y
X0 Y A VP VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 Y A VN VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
.ends

.subckt NAND VP VN A B Y
X0 Y B VP VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X1 VP A Y VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A a_200_10# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=3e+11p ps=2.6e+06u w=1e+06u l=150000u
X3 a_200_10# B VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
.ends


* Top level circuit AND

Xinverter_0 VP VN NAND_0/Y Y inverter
XNAND_0 VP VN A B NAND_0/Y NAND
.end

