* SPICE3 file created from ShiftRegister.ext - technology: sky130A

.subckt inverter A VP VN Y
X0 Y A VN VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
.ends

.subckt DFF D Dn VP VN clk Q Qn
X0 VP a_n390_100# a_n500_n700# VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X1 VN Q Qn VN sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=9.5e+11p ps=5.9e+06u w=1e+06u l=150000u
X2 a_n40_380# Q Qn VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X3 a_n470_n440# a_n390_100# a_n500_n700# VN sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X4 Q Qn a_n40_380# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X5 Qn clk a_n500_n700# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X6 VP clk a_n40_380# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 Q Qn VN VN sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_n390_100# a_n500_n700# a_n470_n440# VN sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X9 Q clk a_n390_100# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X10 a_n500_n700# clk Dn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.5e+11p ps=3.1e+06u w=1e+06u l=600000u
X11 a_n390_100# a_n500_n700# VP VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X12 VN clk a_n470_n440# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 D clk a_n390_100# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=600000u
.ends


* Top level circuit ShiftRegister

Xinverter_0 D VP VN Dn inverter
XDFF_0 D Dn VP VN clk Q3 DFF_1/Dn DFF
XDFF_1 Q3 DFF_1/Dn VP VN clk Q2 DFF_2/Dn DFF
XDFF_2 Q2 DFF_2/Dn VP VN clk Q1 DFF_3/Dn DFF
XDFF_3 Q1 DFF_3/Dn VP VN clk DFF_3/Q Qn0 DFF
.end

