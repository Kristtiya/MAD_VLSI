magic
tech sky130A
timestamp 1614900586
<< nwell >>
rect -275 125 210 440
rect -20 10 210 125
<< nmos >>
rect -200 -65 -185 35
rect -135 -65 -120 35
rect -185 -220 -170 -120
rect -200 -350 -140 -250
rect 50 -185 65 -85
rect 115 -185 130 -85
rect 80 -350 140 -250
<< pmos >>
rect -200 320 -140 420
rect -10 320 50 420
rect -200 145 -185 245
rect -135 145 -120 245
rect 30 190 45 290
rect 55 30 70 130
rect 120 30 135 130
<< ndiff >>
rect -250 20 -200 35
rect -250 -50 -235 20
rect -215 -50 -200 20
rect -250 -65 -200 -50
rect -185 20 -135 35
rect -185 -50 -170 20
rect -150 -50 -135 20
rect -185 -65 -135 -50
rect -120 20 -70 35
rect -120 -50 -105 20
rect -85 -50 -70 20
rect -120 -65 -70 -50
rect -235 -135 -185 -120
rect -235 -205 -220 -135
rect -200 -205 -185 -135
rect -235 -220 -185 -205
rect -170 -135 -120 -120
rect -170 -205 -155 -135
rect -135 -205 -120 -135
rect -170 -220 -120 -205
rect -250 -265 -200 -250
rect -250 -335 -235 -265
rect -215 -335 -200 -265
rect -250 -350 -200 -335
rect -140 -265 -95 -250
rect -140 -335 -130 -265
rect -110 -335 -95 -265
rect -140 -350 -95 -335
rect 0 -100 50 -85
rect 0 -170 15 -100
rect 35 -170 50 -100
rect 0 -185 50 -170
rect 65 -100 115 -85
rect 65 -170 80 -100
rect 100 -170 115 -100
rect 65 -185 115 -170
rect 130 -100 180 -85
rect 130 -170 145 -100
rect 165 -170 180 -100
rect 130 -185 180 -170
rect 30 -265 80 -250
rect 30 -335 45 -265
rect 65 -335 80 -265
rect 30 -350 80 -335
rect 140 -265 190 -250
rect 140 -335 155 -265
rect 175 -335 190 -265
rect 140 -350 190 -335
<< pdiff >>
rect -255 405 -200 420
rect -255 335 -240 405
rect -215 335 -200 405
rect -255 320 -200 335
rect -140 405 -90 420
rect -140 335 -125 405
rect -105 335 -90 405
rect -140 320 -90 335
rect -60 405 -10 420
rect -60 335 -45 405
rect -25 335 -10 405
rect -60 320 -10 335
rect 50 405 100 420
rect 50 335 65 405
rect 85 335 100 405
rect 50 320 100 335
rect -250 230 -200 245
rect -250 160 -235 230
rect -215 160 -200 230
rect -250 145 -200 160
rect -185 230 -135 245
rect -185 160 -170 230
rect -150 160 -135 230
rect -185 145 -135 160
rect -120 230 -70 245
rect -120 160 -105 230
rect -85 160 -70 230
rect -120 145 -70 160
rect -20 275 30 290
rect -20 205 -5 275
rect 15 205 30 275
rect -20 190 30 205
rect 45 275 95 290
rect 45 205 60 275
rect 80 205 95 275
rect 45 190 95 205
rect 5 115 55 130
rect 5 45 20 115
rect 40 45 55 115
rect 5 30 55 45
rect 70 115 120 130
rect 70 45 85 115
rect 105 45 120 115
rect 70 30 120 45
rect 135 115 185 130
rect 135 45 150 115
rect 170 45 185 115
rect 135 30 185 45
<< ndiffc >>
rect -235 -50 -215 20
rect -170 -50 -150 20
rect -105 -50 -85 20
rect -220 -205 -200 -135
rect -155 -205 -135 -135
rect -235 -335 -215 -265
rect -130 -335 -110 -265
rect 15 -170 35 -100
rect 80 -170 100 -100
rect 145 -170 165 -100
rect 45 -335 65 -265
rect 155 -335 175 -265
<< pdiffc >>
rect -240 335 -215 405
rect -125 335 -105 405
rect -45 335 -25 405
rect 65 335 85 405
rect -235 160 -215 230
rect -170 160 -150 230
rect -105 160 -85 230
rect -5 205 15 275
rect 60 205 80 275
rect 20 45 40 115
rect 85 45 105 115
rect 150 45 170 115
<< psubdiff >>
rect -120 -135 -70 -120
rect -120 -205 -105 -135
rect -85 -205 -70 -135
rect -120 -220 -70 -205
<< nsubdiff >>
rect 95 275 145 290
rect 95 205 110 275
rect 130 205 145 275
rect 95 190 145 205
<< psubdiffcont >>
rect -105 -205 -85 -135
<< nsubdiffcont >>
rect 110 205 130 275
<< poly >>
rect -200 420 -140 435
rect -10 420 50 435
rect 155 400 195 410
rect 155 380 165 400
rect 185 380 195 400
rect 155 370 195 380
rect -200 305 -140 320
rect -10 305 50 320
rect -155 300 -140 305
rect -155 285 -35 300
rect 30 290 45 305
rect -200 245 -185 260
rect -135 245 -120 260
rect -50 180 -35 285
rect 30 180 45 190
rect -50 165 45 180
rect 180 175 195 370
rect -200 90 -185 145
rect -135 130 -120 145
rect -160 120 -120 130
rect -160 100 -150 120
rect -130 100 -120 120
rect -160 90 -120 100
rect -225 80 -185 90
rect -225 60 -215 80
rect -195 60 -185 80
rect -225 50 -185 60
rect -200 35 -185 50
rect -135 35 -120 90
rect -200 -80 -185 -65
rect -135 -80 -120 -65
rect -50 -75 -35 165
rect 120 160 195 175
rect 55 130 70 145
rect 120 130 135 160
rect 55 -30 70 30
rect 120 10 135 30
rect 95 0 135 10
rect 95 -20 105 0
rect 125 -20 135 0
rect 95 -30 135 -20
rect 30 -40 70 -30
rect 30 -60 40 -40
rect 60 -60 70 -40
rect 30 -70 70 -60
rect -65 -90 -35 -75
rect 50 -85 65 -70
rect 115 -85 130 -30
rect -185 -120 -170 -105
rect -185 -235 -170 -220
rect -200 -250 -140 -235
rect -200 -365 -140 -350
rect -180 -390 -165 -365
rect -65 -390 -50 -90
rect 50 -200 65 -185
rect 115 -200 130 -185
rect -15 -210 25 -200
rect -15 -230 -5 -210
rect 15 -230 25 -210
rect -15 -240 25 -230
rect -10 -305 5 -240
rect 80 -250 140 -235
rect -25 -315 15 -305
rect -25 -335 -15 -315
rect 5 -335 15 -315
rect -25 -345 15 -335
rect 80 -365 140 -350
rect 80 -390 95 -365
rect -180 -400 -140 -390
rect -180 -420 -170 -400
rect -150 -420 -140 -400
rect -180 -430 -140 -420
rect -80 -400 -40 -390
rect -80 -420 -70 -400
rect -50 -420 -40 -400
rect -80 -430 -40 -420
rect 75 -400 115 -390
rect 75 -420 85 -400
rect 105 -420 115 -400
rect 75 -430 115 -420
<< polycont >>
rect 165 380 185 400
rect -150 100 -130 120
rect -215 60 -195 80
rect 105 -20 125 0
rect 40 -60 60 -40
rect -5 -230 15 -210
rect -15 -335 5 -315
rect -170 -420 -150 -400
rect -70 -420 -50 -400
rect 85 -420 105 -400
<< locali >>
rect -275 445 75 465
rect 55 415 75 445
rect 115 445 210 465
rect -250 410 -205 415
rect -275 405 -205 410
rect -275 390 -240 405
rect -250 335 -240 390
rect -215 335 -205 405
rect -250 325 -205 335
rect -135 405 -95 415
rect -135 335 -125 405
rect -105 335 -95 405
rect -135 325 -95 335
rect -55 405 -15 415
rect -55 335 -45 405
rect -25 335 -15 405
rect -55 325 -15 335
rect 55 405 95 415
rect 55 335 65 405
rect 85 335 95 405
rect 55 325 95 335
rect 115 330 135 445
rect 155 400 210 410
rect 155 380 165 400
rect 185 390 210 400
rect 185 380 195 390
rect 155 370 195 380
rect -135 280 -115 325
rect -55 300 -35 325
rect 115 310 180 330
rect -225 260 -115 280
rect -95 280 -35 300
rect -225 240 -205 260
rect -95 240 -75 280
rect -245 230 -205 240
rect -245 170 -235 230
rect -270 160 -235 170
rect -215 160 -205 230
rect -270 150 -205 160
rect -180 230 -140 240
rect -180 160 -170 230
rect -150 160 -140 230
rect -180 150 -140 160
rect -115 230 -75 240
rect -115 160 -105 230
rect -85 160 -75 230
rect -15 275 25 285
rect -15 205 -5 275
rect 15 205 25 275
rect -15 195 25 205
rect 50 275 140 285
rect 50 205 60 275
rect 80 205 110 275
rect 130 205 140 275
rect 50 195 140 205
rect -115 150 -75 160
rect 5 175 25 195
rect 5 155 110 175
rect -270 130 -250 150
rect -270 120 -120 130
rect -270 110 -150 120
rect -270 30 -250 110
rect -160 100 -150 110
rect -130 100 -120 120
rect -160 90 -120 100
rect -225 80 -185 90
rect -225 60 -215 80
rect -195 70 -185 80
rect -95 70 -75 150
rect 90 125 110 155
rect 160 125 180 310
rect -195 60 -75 70
rect -225 50 -75 60
rect -95 30 -75 50
rect -270 20 -205 30
rect -270 10 -235 20
rect -245 -40 -235 10
rect -270 -50 -235 -40
rect -215 -50 -205 20
rect -270 -60 -205 -50
rect -180 20 -140 30
rect -180 -50 -170 20
rect -150 -50 -140 20
rect -180 -60 -140 -50
rect -115 20 -75 30
rect -115 -50 -105 20
rect -85 -50 -75 20
rect 10 115 50 125
rect 10 45 20 115
rect 40 45 50 115
rect 10 35 50 45
rect 75 115 115 125
rect 75 45 85 115
rect 105 45 115 115
rect 75 35 115 45
rect 140 115 180 125
rect 140 45 150 115
rect 170 45 180 115
rect 140 35 180 45
rect 10 10 30 35
rect -115 -60 -75 -50
rect -270 -255 -250 -60
rect -180 -85 -160 -60
rect -210 -105 -160 -85
rect -95 -85 -75 -60
rect -15 0 135 10
rect -15 -10 105 0
rect -95 -105 -35 -85
rect -210 -125 -190 -105
rect -230 -135 -190 -125
rect -230 -205 -220 -135
rect -200 -205 -190 -135
rect -230 -215 -190 -205
rect -165 -135 -75 -125
rect -165 -205 -155 -135
rect -135 -205 -105 -135
rect -85 -205 -75 -135
rect -165 -215 -75 -205
rect -270 -265 -205 -255
rect -270 -275 -235 -265
rect -245 -335 -235 -275
rect -215 -335 -205 -265
rect -245 -345 -205 -335
rect -135 -265 -100 -255
rect -135 -335 -130 -265
rect -110 -325 -100 -265
rect -55 -265 -35 -105
rect -15 -90 5 -10
rect 95 -20 105 -10
rect 125 -20 135 0
rect 95 -30 135 -20
rect 30 -40 70 -30
rect 30 -60 40 -40
rect 60 -50 70 -40
rect 155 -50 175 35
rect 60 -60 175 -50
rect 30 -70 175 -60
rect 155 -90 175 -70
rect -15 -100 45 -90
rect -15 -110 15 -100
rect 5 -170 15 -110
rect 35 -170 45 -100
rect 5 -180 45 -170
rect 70 -100 110 -90
rect 70 -170 80 -100
rect 100 -170 110 -100
rect 70 -180 110 -170
rect 135 -100 175 -90
rect 135 -170 145 -100
rect 165 -170 175 -100
rect 135 -180 175 -170
rect 5 -200 25 -180
rect -15 -210 25 -200
rect -15 -230 -5 -210
rect 15 -230 25 -210
rect -15 -240 25 -230
rect 145 -255 165 -180
rect 35 -265 75 -255
rect -55 -285 45 -265
rect -25 -315 15 -305
rect -25 -325 -15 -315
rect -110 -335 -15 -325
rect 5 -335 15 -315
rect -135 -345 15 -335
rect 35 -335 45 -285
rect 65 -335 75 -265
rect 35 -345 75 -335
rect 145 -265 185 -255
rect 145 -335 155 -265
rect 175 -335 185 -265
rect 145 -345 185 -335
rect -180 -400 -140 -390
rect -180 -420 -170 -400
rect -150 -420 -140 -400
rect -180 -430 -140 -420
rect -80 -400 -40 -390
rect -80 -420 -70 -400
rect -50 -420 -40 -400
rect -80 -430 -40 -420
rect 75 -400 115 -390
rect 75 -420 85 -400
rect 105 -420 115 -400
rect 75 -430 115 -420
<< viali >>
rect -170 160 -150 230
rect 60 205 80 275
rect 110 205 130 275
rect -155 -205 -135 -135
rect -105 -205 -85 -135
rect 80 -170 100 -100
rect -170 -420 -150 -400
rect -70 -420 -50 -400
rect 85 -420 105 -400
<< metal1 >>
rect -275 275 210 415
rect -275 230 60 275
rect -275 160 -170 230
rect -150 205 60 230
rect 80 205 110 275
rect 130 205 210 275
rect -150 160 210 205
rect -275 150 210 160
rect 10 30 30 45
rect 155 30 175 35
rect -275 -100 210 30
rect -275 -135 80 -100
rect -275 -205 -155 -135
rect -135 -205 -105 -135
rect -85 -170 80 -135
rect 100 -170 210 -100
rect -85 -205 210 -170
rect -275 -345 210 -205
rect -275 -400 210 -390
rect -275 -420 -170 -400
rect -150 -420 -70 -400
rect -50 -420 85 -400
rect 105 -420 210 -400
rect -275 -430 210 -420
<< labels >>
rlabel metal1 -275 -410 -275 -410 7 clk
port 5 w
rlabel metal1 -275 -160 -275 -160 7 VN
port 4 w
rlabel locali -275 455 -275 455 7 D
port 1 w
rlabel metal1 -275 280 -275 280 7 VP
port 3 w
rlabel locali -275 400 -275 400 7 Dn
port 2 w
rlabel locali 210 400 210 400 3 Qn
port 7 e
rlabel locali 210 455 210 455 3 Q
port 6 e
<< end >>
