magic
tech sky130A
timestamp 1614821328
<< nwell >>
rect -275 125 230 605
<< nmos >>
rect -195 -65 -180 35
rect -130 -65 -115 35
rect -130 -220 -115 -120
rect 45 -65 60 35
rect 110 -65 125 35
rect 20 -220 80 -120
rect 20 -350 80 -250
<< pmos >>
rect -155 485 -95 585
rect -200 340 -140 440
rect 60 340 75 440
rect -195 145 -180 245
rect -130 145 -115 245
rect 65 145 80 245
rect 130 145 145 245
<< ndiff >>
rect -245 20 -195 35
rect -245 -50 -230 20
rect -210 -50 -195 20
rect -245 -65 -195 -50
rect -180 20 -130 35
rect -180 -50 -165 20
rect -145 -50 -130 20
rect -180 -65 -130 -50
rect -115 20 -65 35
rect -115 -50 -100 20
rect -80 -50 -65 20
rect -115 -65 -65 -50
rect -180 -135 -130 -120
rect -180 -205 -165 -135
rect -145 -205 -130 -135
rect -180 -220 -130 -205
rect -115 -135 -65 -120
rect -115 -205 -100 -135
rect -80 -205 -65 -135
rect -115 -220 -65 -205
rect -5 20 45 35
rect -5 -50 10 20
rect 30 -50 45 20
rect -5 -65 45 -50
rect 60 20 110 35
rect 60 -50 75 20
rect 95 -50 110 20
rect 60 -65 110 -50
rect 125 20 175 35
rect 125 -50 140 20
rect 160 -50 175 20
rect 125 -65 175 -50
rect -30 -135 20 -120
rect -30 -205 -15 -135
rect 5 -205 20 -135
rect -30 -220 20 -205
rect 80 -135 130 -120
rect 80 -205 95 -135
rect 115 -205 130 -135
rect 80 -220 130 -205
rect -30 -265 20 -250
rect -30 -335 -15 -265
rect 5 -335 20 -265
rect -30 -350 20 -335
rect 80 -265 130 -250
rect 80 -335 95 -265
rect 115 -335 130 -265
rect 80 -350 130 -335
<< pdiff >>
rect -210 570 -155 585
rect -210 500 -195 570
rect -170 500 -155 570
rect -210 485 -155 500
rect -95 570 -45 585
rect -95 500 -80 570
rect -60 500 -45 570
rect -95 485 -45 500
rect -255 425 -200 440
rect -255 355 -240 425
rect -215 355 -200 425
rect -255 340 -200 355
rect -140 425 -90 440
rect -140 355 -125 425
rect -105 355 -90 425
rect -140 340 -90 355
rect 10 425 60 440
rect 10 355 25 425
rect 45 355 60 425
rect 10 340 60 355
rect 75 425 125 440
rect 75 355 90 425
rect 110 355 125 425
rect 75 340 125 355
rect -245 230 -195 245
rect -245 160 -230 230
rect -210 160 -195 230
rect -245 145 -195 160
rect -180 230 -130 245
rect -180 160 -165 230
rect -145 160 -130 230
rect -180 145 -130 160
rect -115 230 -65 245
rect -115 160 -100 230
rect -80 160 -65 230
rect -115 145 -65 160
rect 15 230 65 245
rect 15 160 30 230
rect 50 160 65 230
rect 15 145 65 160
rect 80 230 130 245
rect 80 160 95 230
rect 115 160 130 230
rect 80 145 130 160
rect 145 230 195 245
rect 145 160 160 230
rect 180 160 195 230
rect 145 145 195 160
<< ndiffc >>
rect -230 -50 -210 20
rect -165 -50 -145 20
rect -100 -50 -80 20
rect -165 -205 -145 -135
rect -100 -205 -80 -135
rect 10 -50 30 20
rect 75 -50 95 20
rect 140 -50 160 20
rect -15 -205 5 -135
rect 95 -205 115 -135
rect -15 -335 5 -265
rect 95 -335 115 -265
<< pdiffc >>
rect -195 500 -170 570
rect -80 500 -60 570
rect -240 355 -215 425
rect -125 355 -105 425
rect 25 355 45 425
rect 90 355 110 425
rect -230 160 -210 230
rect -165 160 -145 230
rect -100 160 -80 230
rect 30 160 50 230
rect 95 160 115 230
rect 160 160 180 230
<< psubdiff >>
rect -230 -135 -180 -120
rect -230 -205 -215 -135
rect -195 -205 -180 -135
rect -230 -220 -180 -205
<< nsubdiff >>
rect -40 425 10 440
rect -40 355 -25 425
rect -5 355 10 425
rect -40 340 10 355
<< psubdiffcont >>
rect -215 -205 -195 -135
<< nsubdiffcont >>
rect -25 355 -5 425
<< poly >>
rect -155 585 -95 600
rect -155 470 -95 485
rect -155 455 -140 470
rect -200 440 -140 455
rect 60 440 75 455
rect -200 325 -140 340
rect -155 300 -140 325
rect 60 305 75 340
rect -55 300 75 305
rect -220 290 -180 300
rect -220 270 -210 290
rect -190 270 -180 290
rect -155 285 75 300
rect 130 295 230 305
rect 130 290 200 295
rect -220 260 -180 270
rect -195 245 -180 260
rect -130 245 -115 260
rect -195 90 -180 145
rect -130 130 -115 145
rect -155 120 -115 130
rect -155 100 -145 120
rect -125 100 -115 120
rect -155 90 -115 100
rect -220 80 -180 90
rect -220 60 -210 80
rect -190 60 -180 80
rect -220 50 -180 60
rect -195 35 -180 50
rect -130 35 -115 90
rect -195 -80 -180 -65
rect -130 -80 -115 -65
rect -130 -120 -115 -105
rect -130 -235 -115 -220
rect -55 -235 -40 285
rect 65 245 80 260
rect 130 245 145 290
rect 190 275 200 290
rect 220 275 230 295
rect 190 265 230 275
rect 65 130 80 145
rect 130 130 145 145
rect 45 115 80 130
rect 110 120 150 130
rect 45 90 60 115
rect 110 100 120 120
rect 140 100 150 120
rect 110 90 150 100
rect 45 80 85 90
rect 45 60 55 80
rect 75 60 85 80
rect 45 50 85 60
rect 45 35 60 50
rect 110 35 125 90
rect 45 -80 60 -65
rect 110 -80 125 -65
rect 110 -95 160 -80
rect 20 -120 80 -105
rect -130 -250 -40 -235
rect 20 -250 80 -220
rect -130 -390 -115 -250
rect 145 -255 160 -95
rect 145 -265 185 -255
rect 145 -285 155 -265
rect 175 -285 185 -265
rect 145 -295 185 -285
rect 20 -365 80 -350
rect 40 -390 55 -365
rect -155 -400 -115 -390
rect -155 -420 -145 -400
rect -125 -420 -115 -400
rect -155 -430 -115 -420
rect 15 -400 55 -390
rect 15 -420 25 -400
rect 45 -420 55 -400
rect 15 -430 55 -420
<< polycont >>
rect -210 270 -190 290
rect -145 100 -125 120
rect -210 60 -190 80
rect 200 275 220 295
rect 120 100 140 120
rect 55 60 75 80
rect 155 -285 175 -265
rect -145 -420 -125 -400
rect 25 -420 45 -400
<< locali >>
rect -275 650 -185 670
rect -275 610 -230 630
rect -250 435 -230 610
rect -205 580 -185 650
rect 150 650 230 670
rect -205 570 -160 580
rect -205 500 -195 570
rect -170 500 -160 570
rect -205 490 -160 500
rect -90 570 -50 580
rect -90 500 -80 570
rect -60 500 -50 570
rect -90 490 -50 500
rect -250 425 -205 435
rect -250 355 -240 425
rect -215 355 -205 425
rect -250 345 -205 355
rect -135 425 -95 435
rect -135 355 -125 425
rect -105 355 -95 425
rect -135 345 -95 355
rect -130 325 -110 345
rect -75 325 -55 490
rect -35 425 55 435
rect -35 355 -25 425
rect -5 355 25 425
rect 45 355 55 425
rect -35 345 55 355
rect 80 425 120 435
rect 80 355 90 425
rect 110 355 120 425
rect 80 345 120 355
rect -200 305 -110 325
rect -90 305 -55 325
rect -200 300 -180 305
rect -220 290 -180 300
rect -220 270 -210 290
rect -190 270 -180 290
rect -220 260 -180 270
rect -90 240 -70 305
rect 85 240 105 345
rect 150 240 170 650
rect 190 610 230 630
rect 190 305 210 610
rect 190 295 230 305
rect 190 275 200 295
rect 220 275 230 295
rect 190 265 230 275
rect -240 230 -200 240
rect -240 170 -230 230
rect -270 160 -230 170
rect -210 160 -200 230
rect -270 150 -200 160
rect -175 230 -135 240
rect -175 160 -165 230
rect -145 160 -135 230
rect -175 150 -135 160
rect -110 230 -70 240
rect -110 160 -100 230
rect -80 160 -70 230
rect -110 150 -70 160
rect -270 130 -250 150
rect -270 120 -115 130
rect -270 110 -145 120
rect -270 30 -250 110
rect -155 100 -145 110
rect -125 100 -115 120
rect -155 90 -115 100
rect -220 80 -180 90
rect -220 60 -210 80
rect -190 70 -180 80
rect -90 70 -70 150
rect 20 230 60 240
rect 20 160 30 230
rect 50 160 60 230
rect 20 150 60 160
rect 85 230 125 240
rect 85 160 95 230
rect 115 160 125 230
rect 85 150 125 160
rect 150 230 190 240
rect 150 160 160 230
rect 180 160 190 230
rect 150 150 190 160
rect 20 130 40 150
rect 0 120 150 130
rect 0 110 120 120
rect -190 60 -20 70
rect -220 50 -20 60
rect -90 30 -70 50
rect -270 20 -200 30
rect -270 10 -230 20
rect -240 -40 -230 10
rect -270 -50 -230 -40
rect -210 -50 -200 20
rect -270 -60 -200 -50
rect -175 20 -135 30
rect -175 -50 -165 20
rect -145 -50 -135 20
rect -175 -60 -135 -50
rect -110 20 -70 30
rect -110 -50 -100 20
rect -80 -50 -70 20
rect -110 -60 -70 -50
rect -270 -255 -250 -60
rect -155 -80 -135 -60
rect -155 -100 -90 -80
rect -110 -125 -90 -100
rect -40 -90 -20 50
rect 0 30 20 110
rect 110 100 120 110
rect 140 100 150 120
rect 110 90 150 100
rect 45 80 85 90
rect 45 60 55 80
rect 75 70 85 80
rect 170 70 190 150
rect 75 60 210 70
rect 45 50 210 60
rect 150 30 170 50
rect 0 20 40 30
rect 0 -50 10 20
rect 30 -50 40 20
rect 0 -60 40 -50
rect 65 20 105 30
rect 65 -50 75 20
rect 95 -50 105 20
rect 65 -60 105 -50
rect 130 20 170 30
rect 130 -50 140 20
rect 160 -50 170 20
rect 130 -60 170 -50
rect -40 -110 -5 -90
rect -25 -125 -5 -110
rect 190 -125 210 50
rect -225 -135 -135 -125
rect -225 -205 -215 -135
rect -195 -205 -165 -135
rect -145 -205 -135 -135
rect -225 -215 -135 -205
rect -110 -135 -70 -125
rect -110 -205 -100 -135
rect -80 -205 -70 -135
rect -110 -215 -70 -205
rect -25 -135 15 -125
rect -25 -205 -15 -135
rect 5 -205 15 -135
rect -25 -215 15 -205
rect 85 -135 210 -125
rect 85 -205 95 -135
rect 115 -145 210 -135
rect 115 -205 125 -145
rect 85 -215 125 -205
rect -270 -265 15 -255
rect -270 -275 -15 -265
rect -25 -335 -15 -275
rect 5 -335 15 -265
rect -25 -345 15 -335
rect 85 -265 185 -255
rect 85 -335 95 -265
rect 115 -275 155 -265
rect 115 -335 125 -275
rect 145 -285 155 -275
rect 175 -285 185 -265
rect 145 -295 185 -285
rect 85 -345 125 -335
rect -155 -400 -115 -390
rect -155 -420 -145 -400
rect -125 -420 -115 -400
rect -155 -430 -115 -420
rect 15 -400 55 -390
rect 15 -420 25 -400
rect 45 -420 55 -400
rect 15 -430 55 -420
<< viali >>
rect -25 355 -5 425
rect 25 355 45 425
rect -165 160 -145 230
rect 75 -50 95 20
rect -215 -205 -195 -135
rect -165 -205 -145 -135
<< metal1 >>
rect -275 425 230 580
rect -275 355 -25 425
rect -5 355 25 425
rect 45 355 230 425
rect -275 230 230 355
rect -275 160 -165 230
rect -145 160 230 230
rect -275 150 230 160
rect -275 20 230 30
rect -275 -50 75 20
rect 95 -50 230 20
rect -275 -135 230 -50
rect -275 -205 -215 -135
rect -195 -205 -165 -135
rect -145 -205 230 -135
rect -275 -345 230 -205
rect -275 -430 230 -390
<< labels >>
rlabel metal1 -275 370 -275 370 7 VP
port 4 w
rlabel metal1 -275 -160 -275 -160 3 VN
port 5 e
rlabel metal1 -275 -410 -275 -410 7 clk
port 3 w
rlabel locali -275 660 -275 660 7 D
port 1 w
rlabel locali -275 620 -275 620 7 Dn
port 2 w
rlabel locali 230 660 230 660 3 Q
port 6 e
rlabel locali 230 620 230 620 3 Qn
port 7 e
<< end >>
