magic
tech sky130A
timestamp 1614901737
<< nwell >>
rect 280 570 485 835
<< nmos >>
rect 400 335 415 435
<< pmos >>
rect 400 590 415 690
<< ndiff >>
rect 350 420 400 435
rect 350 350 365 420
rect 385 350 400 420
rect 350 335 400 350
rect 415 420 465 435
rect 415 350 430 420
rect 450 350 465 420
rect 415 335 465 350
<< pdiff >>
rect 350 675 400 690
rect 350 605 365 675
rect 385 605 400 675
rect 350 590 400 605
rect 415 675 465 690
rect 415 605 430 675
rect 450 605 465 675
rect 415 590 465 605
<< ndiffc >>
rect 365 350 385 420
rect 430 350 450 420
<< pdiffc >>
rect 365 605 385 675
rect 430 605 450 675
<< psubdiff >>
rect 300 420 350 435
rect 300 350 315 420
rect 335 350 350 420
rect 300 335 350 350
<< nsubdiff >>
rect 300 675 350 690
rect 300 605 315 675
rect 335 605 350 675
rect 300 590 350 605
<< psubdiffcont >>
rect 315 350 335 420
<< nsubdiffcont >>
rect 315 605 335 675
<< poly >>
rect 380 735 420 745
rect 380 715 390 735
rect 410 715 420 735
rect 380 705 420 715
rect 400 690 415 705
rect 400 435 415 590
rect 400 320 415 335
<< polycont >>
rect 390 715 410 735
<< locali >>
rect 400 865 485 885
rect 400 745 420 865
rect 380 735 420 745
rect 380 725 390 735
rect 280 715 390 725
rect 410 715 420 735
rect 280 705 420 715
rect 440 810 485 830
rect 440 685 460 810
rect 305 675 395 685
rect 305 605 315 675
rect 335 605 365 675
rect 385 605 395 675
rect 305 595 395 605
rect 420 675 460 685
rect 420 605 430 675
rect 450 605 460 675
rect 420 595 460 605
rect 440 430 460 595
rect 305 420 395 430
rect 305 350 315 420
rect 335 350 365 420
rect 385 350 395 420
rect 305 340 395 350
rect 420 420 460 430
rect 420 350 430 420
rect 450 350 460 420
rect 420 340 460 350
<< viali >>
rect 315 605 335 675
rect 365 605 385 675
rect 315 350 335 420
rect 365 350 385 420
<< metal1 >>
rect 280 675 485 835
rect 280 605 315 675
rect 335 605 365 675
rect 385 605 485 675
rect 280 570 485 605
rect 280 420 485 450
rect 280 350 315 420
rect 335 350 365 420
rect 385 350 485 420
rect 280 75 485 350
<< labels >>
rlabel locali 280 715 280 715 7 A
port 1 w
rlabel metal1 280 700 280 700 7 VP
port 2 w
rlabel metal1 280 270 280 270 7 VN
port 3 w
rlabel locali 485 820 485 820 3 Y
port 4 e
<< end >>
