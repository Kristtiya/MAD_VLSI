magic
tech sky130A
timestamp 1618101028
<< nwell >>
rect 1210 -150 3265 1090
rect 2990 -1650 3265 -150
<< nmos >>
rect 1295 -1630 1345 -430
rect 1395 -1630 1445 -430
rect 1495 -1630 1545 -430
rect 1595 -1630 1645 -430
rect 1695 -1630 1745 -430
rect 1795 -1630 1845 -430
rect 1995 -1630 2045 -430
rect 2095 -1630 2145 -430
rect 2195 -1630 2245 -430
rect 2295 -1630 2345 -430
rect 2395 -1630 2445 -430
rect 2625 -1630 2675 -430
rect 2855 -1630 2905 -430
<< pmos >>
rect 1330 -130 1380 1070
rect 1430 -130 1480 1070
rect 1530 -130 1580 1070
rect 1630 -130 1680 1070
rect 1730 -130 1780 1070
rect 1830 -130 1880 1070
rect 1930 -130 1980 1070
rect 2130 -130 2180 1070
rect 2230 -130 2280 1070
rect 2330 -130 2380 1070
rect 2430 -130 2480 1070
rect 2530 -130 2580 1070
rect 2630 -130 2680 1070
rect 2730 -130 2780 1070
rect 2960 -130 3010 1070
rect 3060 -130 3110 1070
rect 3060 -1630 3110 -430
<< ndiff >>
rect 1245 -445 1295 -430
rect 1245 -1615 1260 -445
rect 1280 -1615 1295 -445
rect 1245 -1630 1295 -1615
rect 1345 -445 1395 -430
rect 1345 -1615 1360 -445
rect 1380 -1615 1395 -445
rect 1345 -1630 1395 -1615
rect 1445 -445 1495 -430
rect 1445 -1615 1460 -445
rect 1480 -1615 1495 -445
rect 1445 -1630 1495 -1615
rect 1545 -445 1595 -430
rect 1545 -1615 1560 -445
rect 1580 -1615 1595 -445
rect 1545 -1630 1595 -1615
rect 1645 -445 1695 -430
rect 1645 -1615 1660 -445
rect 1680 -1615 1695 -445
rect 1645 -1630 1695 -1615
rect 1745 -445 1795 -430
rect 1745 -1615 1760 -445
rect 1780 -1615 1795 -445
rect 1745 -1630 1795 -1615
rect 1845 -445 1895 -430
rect 1945 -445 1995 -430
rect 1845 -1615 1860 -445
rect 1880 -1615 1895 -445
rect 1945 -1615 1960 -445
rect 1980 -1615 1995 -445
rect 1845 -1630 1895 -1615
rect 1945 -1630 1995 -1615
rect 2045 -445 2095 -430
rect 2045 -1615 2060 -445
rect 2080 -1615 2095 -445
rect 2045 -1630 2095 -1615
rect 2145 -445 2195 -430
rect 2145 -1615 2160 -445
rect 2180 -1615 2195 -445
rect 2145 -1630 2195 -1615
rect 2245 -445 2295 -430
rect 2245 -1615 2260 -445
rect 2280 -1615 2295 -445
rect 2245 -1630 2295 -1615
rect 2345 -445 2395 -430
rect 2345 -1615 2360 -445
rect 2380 -1615 2395 -445
rect 2345 -1630 2395 -1615
rect 2445 -445 2495 -430
rect 2445 -1615 2460 -445
rect 2480 -1615 2495 -445
rect 2445 -1630 2495 -1615
rect 2575 -445 2625 -430
rect 2575 -1615 2590 -445
rect 2610 -1615 2625 -445
rect 2575 -1630 2625 -1615
rect 2675 -445 2725 -430
rect 2675 -1615 2690 -445
rect 2710 -1615 2725 -445
rect 2675 -1630 2725 -1615
rect 2805 -445 2855 -430
rect 2805 -1615 2820 -445
rect 2840 -1615 2855 -445
rect 2805 -1630 2855 -1615
rect 2905 -445 2955 -430
rect 2905 -1615 2920 -445
rect 2940 -1615 2955 -445
rect 2905 -1630 2955 -1615
<< pdiff >>
rect 1280 1055 1330 1070
rect 1280 -115 1295 1055
rect 1315 -115 1330 1055
rect 1280 -130 1330 -115
rect 1380 1055 1430 1070
rect 1380 -115 1395 1055
rect 1415 -115 1430 1055
rect 1380 -130 1430 -115
rect 1480 1055 1530 1070
rect 1480 -115 1495 1055
rect 1515 -115 1530 1055
rect 1480 -130 1530 -115
rect 1580 1055 1630 1070
rect 1580 -115 1595 1055
rect 1615 -115 1630 1055
rect 1580 -130 1630 -115
rect 1680 1055 1730 1070
rect 1680 -115 1695 1055
rect 1715 -115 1730 1055
rect 1680 -130 1730 -115
rect 1780 1055 1830 1070
rect 1780 -115 1795 1055
rect 1815 -115 1830 1055
rect 1780 -130 1830 -115
rect 1880 1055 1930 1070
rect 1880 -115 1895 1055
rect 1915 -115 1930 1055
rect 1880 -130 1930 -115
rect 1980 1055 2030 1070
rect 2080 1055 2130 1070
rect 1980 -115 1995 1055
rect 2015 -115 2030 1055
rect 2080 -115 2095 1055
rect 2115 -115 2130 1055
rect 1980 -130 2030 -115
rect 2080 -130 2130 -115
rect 2180 1055 2230 1070
rect 2180 -115 2195 1055
rect 2215 -115 2230 1055
rect 2180 -130 2230 -115
rect 2280 1055 2330 1070
rect 2280 -115 2295 1055
rect 2315 -115 2330 1055
rect 2280 -130 2330 -115
rect 2380 1055 2430 1070
rect 2380 -115 2395 1055
rect 2415 -115 2430 1055
rect 2380 -130 2430 -115
rect 2480 1055 2530 1070
rect 2480 -115 2495 1055
rect 2515 -115 2530 1055
rect 2480 -130 2530 -115
rect 2580 1055 2630 1070
rect 2580 -115 2595 1055
rect 2615 -115 2630 1055
rect 2580 -130 2630 -115
rect 2680 1055 2730 1070
rect 2680 -115 2695 1055
rect 2715 -115 2730 1055
rect 2680 -130 2730 -115
rect 2780 1055 2830 1070
rect 2780 -115 2795 1055
rect 2815 -115 2830 1055
rect 2780 -130 2830 -115
rect 2910 1055 2960 1070
rect 2910 -115 2925 1055
rect 2945 -115 2960 1055
rect 2910 -130 2960 -115
rect 3010 1055 3060 1070
rect 3010 -115 3025 1055
rect 3045 -115 3060 1055
rect 3010 -130 3060 -115
rect 3110 1055 3160 1070
rect 3110 -115 3125 1055
rect 3145 -115 3160 1055
rect 3110 -130 3160 -115
rect 3010 -445 3060 -430
rect 3010 -1615 3025 -445
rect 3045 -1615 3060 -445
rect 3010 -1630 3060 -1615
rect 3110 -445 3160 -430
rect 3110 -1615 3125 -445
rect 3145 -1615 3160 -445
rect 3110 -1630 3160 -1615
<< ndiffc >>
rect 1260 -1615 1280 -445
rect 1360 -1615 1380 -445
rect 1460 -1615 1480 -445
rect 1560 -1615 1580 -445
rect 1660 -1615 1680 -445
rect 1760 -1615 1780 -445
rect 1860 -1615 1880 -445
rect 1960 -1615 1980 -445
rect 2060 -1615 2080 -445
rect 2160 -1615 2180 -445
rect 2260 -1615 2280 -445
rect 2360 -1615 2380 -445
rect 2460 -1615 2480 -445
rect 2590 -1615 2610 -445
rect 2690 -1615 2710 -445
rect 2820 -1615 2840 -445
rect 2920 -1615 2940 -445
<< pdiffc >>
rect 1295 -115 1315 1055
rect 1395 -115 1415 1055
rect 1495 -115 1515 1055
rect 1595 -115 1615 1055
rect 1695 -115 1715 1055
rect 1795 -115 1815 1055
rect 1895 -115 1915 1055
rect 1995 -115 2015 1055
rect 2095 -115 2115 1055
rect 2195 -115 2215 1055
rect 2295 -115 2315 1055
rect 2395 -115 2415 1055
rect 2495 -115 2515 1055
rect 2595 -115 2615 1055
rect 2695 -115 2715 1055
rect 2795 -115 2815 1055
rect 2925 -115 2945 1055
rect 3025 -115 3045 1055
rect 3125 -115 3145 1055
rect 3025 -1615 3045 -445
rect 3125 -1615 3145 -445
<< psubdiff >>
rect 1895 -445 1945 -430
rect 1895 -1615 1910 -445
rect 1930 -1615 1945 -445
rect 1895 -1630 1945 -1615
rect 2525 -445 2575 -430
rect 2525 -1615 2540 -445
rect 2560 -1615 2575 -445
rect 2525 -1630 2575 -1615
rect 2755 -445 2805 -430
rect 2755 -1615 2770 -445
rect 2790 -1615 2805 -445
rect 2755 -1630 2805 -1615
<< nsubdiff >>
rect 1230 1055 1280 1070
rect 1230 -115 1245 1055
rect 1265 -115 1280 1055
rect 1230 -130 1280 -115
rect 2030 1055 2080 1070
rect 2030 -115 2045 1055
rect 2065 -115 2080 1055
rect 2030 -130 2080 -115
rect 2830 1055 2880 1070
rect 2830 -115 2845 1055
rect 2865 -115 2880 1055
rect 2830 -130 2880 -115
rect 3160 -445 3210 -430
rect 3160 -1615 3175 -445
rect 3195 -1615 3210 -445
rect 3160 -1630 3210 -1615
<< psubdiffcont >>
rect 1910 -1615 1930 -445
rect 2540 -1615 2560 -445
rect 2770 -1615 2790 -445
<< nsubdiffcont >>
rect 1245 -115 1265 1055
rect 2045 -115 2065 1055
rect 2845 -115 2865 1055
rect 3175 -1615 3195 -445
<< poly >>
rect 1830 1150 2280 1165
rect 1285 1115 1325 1125
rect 1285 1095 1295 1115
rect 1315 1100 1325 1115
rect 1830 1100 1880 1150
rect 2035 1115 2075 1125
rect 2035 1100 2045 1115
rect 1315 1095 1380 1100
rect 1285 1085 1380 1095
rect 1330 1070 1380 1085
rect 1430 1085 1880 1100
rect 1430 1070 1480 1085
rect 1530 1070 1580 1085
rect 1630 1070 1680 1085
rect 1730 1070 1780 1085
rect 1830 1070 1880 1085
rect 1930 1095 2045 1100
rect 2065 1100 2075 1115
rect 2230 1100 2280 1150
rect 2785 1115 2825 1125
rect 2785 1100 2795 1115
rect 2065 1095 2180 1100
rect 1930 1085 2180 1095
rect 1930 1070 1980 1085
rect 2130 1070 2180 1085
rect 2230 1085 2680 1100
rect 2230 1070 2280 1085
rect 2330 1070 2380 1085
rect 2430 1070 2480 1085
rect 2530 1070 2580 1085
rect 2630 1070 2680 1085
rect 2730 1095 2795 1100
rect 2815 1095 2825 1115
rect 2730 1085 2825 1095
rect 2960 1085 3110 1105
rect 2730 1070 2780 1085
rect 2960 1070 3010 1085
rect 3060 1070 3110 1085
rect 3185 -110 3225 -100
rect 3185 -130 3195 -110
rect 3215 -130 3225 -110
rect 1330 -145 1380 -130
rect 1430 -145 1480 -130
rect 1530 -145 1580 -130
rect 1630 -155 1680 -130
rect 1730 -145 1780 -130
rect 1830 -145 1880 -130
rect 1930 -145 1980 -130
rect 2130 -145 2180 -130
rect 2230 -145 2280 -130
rect 2330 -145 2380 -130
rect 2430 -145 2480 -130
rect 2530 -145 2580 -130
rect 2630 -145 2680 -130
rect 2730 -145 2780 -130
rect 2960 -145 3010 -130
rect 3060 -145 3110 -130
rect 3185 -140 3225 -130
rect 1630 -185 1640 -155
rect 1670 -185 1680 -155
rect 1630 -195 1680 -185
rect 2005 -160 2045 -150
rect 2005 -180 2015 -160
rect 2035 -170 2045 -160
rect 2035 -180 2345 -170
rect 2005 -185 2315 -180
rect 2005 -190 2045 -185
rect 1645 -235 1660 -195
rect 2305 -200 2315 -185
rect 2335 -200 2345 -180
rect 3065 -180 3105 -170
rect 3065 -195 3075 -180
rect 2305 -210 2345 -200
rect 2380 -200 3075 -195
rect 3095 -200 3105 -180
rect 2380 -210 3105 -200
rect 2380 -235 2395 -210
rect 1645 -250 2395 -235
rect 2855 -245 3105 -235
rect 2855 -250 3075 -245
rect 2295 -375 2345 -365
rect 1900 -385 1940 -375
rect 1900 -400 1910 -385
rect 1795 -405 1910 -400
rect 1930 -400 1940 -385
rect 2150 -385 2190 -375
rect 2150 -400 2160 -385
rect 1930 -405 2045 -400
rect 1795 -415 2045 -405
rect 1295 -430 1345 -415
rect 1395 -430 1445 -415
rect 1495 -430 1545 -415
rect 1595 -430 1645 -415
rect 1695 -430 1745 -415
rect 1795 -430 1845 -415
rect 1995 -430 2045 -415
rect 2095 -405 2160 -400
rect 2180 -400 2190 -385
rect 2180 -405 2245 -400
rect 2095 -415 2245 -405
rect 2095 -430 2145 -415
rect 2195 -430 2245 -415
rect 2295 -405 2305 -375
rect 2335 -405 2345 -375
rect 2295 -430 2345 -405
rect 2395 -375 2445 -365
rect 2395 -405 2405 -375
rect 2435 -405 2445 -375
rect 2395 -430 2445 -405
rect 2530 -385 2570 -375
rect 2530 -405 2540 -385
rect 2560 -400 2570 -385
rect 2560 -405 2675 -400
rect 2530 -415 2675 -405
rect 2625 -430 2675 -415
rect 2855 -415 2870 -250
rect 3065 -265 3075 -250
rect 3095 -265 3105 -245
rect 3065 -275 3105 -265
rect 2930 -285 2970 -275
rect 2930 -305 2940 -285
rect 2960 -305 2970 -285
rect 2930 -315 2970 -305
rect 2995 -285 3035 -275
rect 2995 -305 3005 -285
rect 3025 -305 3035 -285
rect 2995 -315 3035 -305
rect 2930 -375 2945 -315
rect 2995 -375 3010 -315
rect 2930 -385 2970 -375
rect 2930 -405 2940 -385
rect 2960 -405 2970 -385
rect 2930 -415 2970 -405
rect 2995 -385 3035 -375
rect 2995 -405 3005 -385
rect 3025 -405 3035 -385
rect 2995 -415 3035 -405
rect 3185 -380 3200 -140
rect 3185 -390 3225 -380
rect 3185 -410 3195 -390
rect 3215 -410 3225 -390
rect 2855 -430 2905 -415
rect 3060 -430 3110 -415
rect 3185 -420 3225 -410
rect 1295 -1645 1345 -1630
rect 1250 -1655 1345 -1645
rect 1250 -1675 1260 -1655
rect 1280 -1660 1345 -1655
rect 1280 -1675 1290 -1660
rect 1250 -1685 1290 -1675
rect 1395 -1670 1445 -1630
rect 1495 -1670 1545 -1630
rect 1595 -1670 1645 -1630
rect 1695 -1670 1745 -1630
rect 1795 -1645 1845 -1630
rect 1995 -1645 2045 -1630
rect 2095 -1645 2145 -1630
rect 2195 -1645 2245 -1630
rect 2295 -1670 2345 -1630
rect 2395 -1645 2445 -1630
rect 2625 -1645 2675 -1630
rect 2855 -1670 2905 -1630
rect 1395 -1685 2905 -1670
rect 3060 -1665 3110 -1630
rect 3060 -1695 3070 -1665
rect 3100 -1695 3110 -1665
rect 3060 -1705 3110 -1695
<< polycont >>
rect 1295 1095 1315 1115
rect 2045 1095 2065 1115
rect 2795 1095 2815 1115
rect 3195 -130 3215 -110
rect 1640 -185 1670 -155
rect 2015 -180 2035 -160
rect 2315 -200 2335 -180
rect 3075 -200 3095 -180
rect 1910 -405 1930 -385
rect 2160 -405 2180 -385
rect 2305 -405 2335 -375
rect 2405 -405 2435 -375
rect 2540 -405 2560 -385
rect 3075 -265 3095 -245
rect 2940 -305 2960 -285
rect 3005 -305 3025 -285
rect 2940 -405 2960 -385
rect 3005 -405 3025 -385
rect 3195 -410 3215 -390
rect 1260 -1675 1280 -1655
rect 3070 -1695 3100 -1665
<< locali >>
rect 1390 1135 1820 1165
rect 1285 1115 1325 1125
rect 1285 1095 1295 1115
rect 1315 1095 1325 1115
rect 1285 1065 1325 1095
rect 1390 1065 1420 1135
rect 1590 1065 1620 1135
rect 1790 1065 1820 1135
rect 2035 1115 2075 1125
rect 2035 1095 2045 1115
rect 2065 1095 2075 1115
rect 2035 1065 2075 1095
rect 2295 1100 2715 1120
rect 2295 1065 2315 1100
rect 2495 1065 2515 1100
rect 2695 1065 2715 1100
rect 2785 1115 2825 1125
rect 2785 1095 2795 1115
rect 2815 1095 2825 1115
rect 2785 1085 2825 1095
rect 2785 1065 2820 1085
rect 1235 1055 1325 1065
rect 1235 -115 1245 1055
rect 1265 -115 1295 1055
rect 1315 -115 1325 1055
rect 1235 -125 1325 -115
rect 1385 1055 1425 1065
rect 1385 -115 1395 1055
rect 1415 -115 1425 1055
rect 1385 -125 1425 -115
rect 1485 1055 1525 1065
rect 1485 -115 1495 1055
rect 1515 -115 1525 1055
rect 1485 -125 1525 -115
rect 1585 1055 1625 1065
rect 1585 -115 1595 1055
rect 1615 -115 1625 1055
rect 1585 -125 1625 -115
rect 1685 1055 1725 1065
rect 1685 -115 1695 1055
rect 1715 -115 1725 1055
rect 1685 -125 1725 -115
rect 1785 1055 1825 1065
rect 1785 -115 1795 1055
rect 1815 -115 1825 1055
rect 1785 -125 1825 -115
rect 1885 1055 1925 1065
rect 1885 -115 1895 1055
rect 1915 -115 1925 1055
rect 1885 -125 1925 -115
rect 1985 1055 2125 1065
rect 1985 -115 1995 1055
rect 2015 -115 2045 1055
rect 2065 -115 2095 1055
rect 2115 -115 2125 1055
rect 1985 -125 2125 -115
rect 2185 1055 2225 1065
rect 2185 -115 2195 1055
rect 2215 -115 2225 1055
rect 2185 -125 2225 -115
rect 2285 1055 2325 1065
rect 2285 -115 2295 1055
rect 2315 -115 2325 1055
rect 2285 -125 2325 -115
rect 2385 1055 2425 1065
rect 2385 -115 2395 1055
rect 2415 -115 2425 1055
rect 2385 -125 2425 -115
rect 2485 1055 2525 1065
rect 2485 -115 2495 1055
rect 2515 -115 2525 1055
rect 2485 -125 2525 -115
rect 2585 1055 2625 1065
rect 2585 -115 2595 1055
rect 2615 -115 2625 1055
rect 2585 -125 2625 -115
rect 2685 1055 2725 1065
rect 2685 -115 2695 1055
rect 2715 -115 2725 1055
rect 2685 -125 2725 -115
rect 2785 1055 2875 1065
rect 2785 -115 2795 1055
rect 2815 -115 2845 1055
rect 2865 -115 2875 1055
rect 2785 -125 2875 -115
rect 2915 1055 2955 1065
rect 2915 -115 2925 1055
rect 2945 -115 2955 1055
rect 2915 -125 2955 -115
rect 3015 1055 3055 1065
rect 3015 -115 3025 1055
rect 3045 -115 3055 1055
rect 3015 -125 3055 -115
rect 3115 1055 3155 1065
rect 3115 -115 3125 1055
rect 3145 -115 3155 1055
rect 3115 -125 3155 -115
rect 3185 -105 3225 -100
rect 3185 -110 3265 -105
rect 1495 -145 1515 -125
rect 1695 -145 1715 -125
rect 1210 -155 1715 -145
rect 1210 -165 1640 -155
rect 1630 -185 1640 -165
rect 1670 -165 1715 -155
rect 1895 -150 1915 -125
rect 2195 -145 2215 -125
rect 1895 -160 2045 -150
rect 1670 -185 1680 -165
rect 1895 -170 2015 -160
rect 1630 -195 1680 -185
rect 2005 -180 2015 -170
rect 2035 -180 2045 -160
rect 2005 -190 2045 -180
rect 2160 -165 2215 -145
rect 2395 -145 2415 -125
rect 2595 -145 2615 -125
rect 2395 -165 2615 -145
rect 2160 -375 2180 -165
rect 2305 -180 2345 -170
rect 2305 -200 2315 -180
rect 2335 -200 2345 -180
rect 2305 -210 2345 -200
rect 2315 -365 2335 -210
rect 2295 -375 2345 -365
rect 1900 -385 1940 -375
rect 1360 -415 1780 -395
rect 1360 -435 1380 -415
rect 1560 -435 1580 -415
rect 1760 -435 1780 -415
rect 1900 -405 1910 -385
rect 1930 -405 1940 -385
rect 1900 -435 1940 -405
rect 2070 -385 2190 -375
rect 2070 -400 2160 -385
rect 2070 -435 2090 -400
rect 2150 -405 2160 -400
rect 2180 -405 2190 -385
rect 2150 -415 2190 -405
rect 2295 -405 2305 -375
rect 2335 -395 2345 -375
rect 2395 -375 2445 -365
rect 2335 -405 2370 -395
rect 2295 -415 2370 -405
rect 2395 -405 2405 -375
rect 2435 -395 2445 -375
rect 2530 -375 2550 -165
rect 2930 -275 2950 -125
rect 3015 -275 3035 -125
rect 3185 -130 3195 -110
rect 3215 -125 3265 -110
rect 3215 -130 3225 -125
rect 3185 -140 3225 -130
rect 3065 -180 3265 -170
rect 3065 -200 3075 -180
rect 3095 -190 3265 -180
rect 3095 -200 3105 -190
rect 3065 -210 3105 -200
rect 3065 -245 3265 -235
rect 3065 -265 3075 -245
rect 3095 -255 3265 -245
rect 3095 -265 3105 -255
rect 3065 -275 3105 -265
rect 2930 -285 2970 -275
rect 2930 -305 2940 -285
rect 2960 -305 2970 -285
rect 2930 -315 2970 -305
rect 2995 -285 3035 -275
rect 2995 -305 3005 -285
rect 3025 -305 3035 -285
rect 2995 -315 3035 -305
rect 3115 -320 3265 -300
rect 3115 -335 3135 -320
rect 2835 -355 3135 -335
rect 2530 -380 2570 -375
rect 2835 -380 2855 -355
rect 2530 -385 2855 -380
rect 2435 -405 2470 -395
rect 2395 -415 2470 -405
rect 2350 -435 2370 -415
rect 2450 -435 2470 -415
rect 2530 -405 2540 -385
rect 2560 -400 2855 -385
rect 2930 -385 2970 -375
rect 2560 -405 2570 -400
rect 2530 -435 2570 -405
rect 2930 -405 2940 -385
rect 2960 -405 2970 -385
rect 2930 -415 2970 -405
rect 2995 -385 3035 -375
rect 2995 -405 3005 -385
rect 3025 -405 3035 -385
rect 2995 -415 3035 -405
rect 2930 -435 2950 -415
rect 1250 -445 1290 -435
rect 1250 -1615 1260 -445
rect 1280 -1615 1290 -445
rect 1250 -1655 1290 -1615
rect 1350 -445 1390 -435
rect 1350 -1615 1360 -445
rect 1380 -1615 1390 -445
rect 1350 -1625 1390 -1615
rect 1450 -445 1490 -435
rect 1450 -1615 1460 -445
rect 1480 -1615 1490 -445
rect 1450 -1625 1490 -1615
rect 1550 -445 1590 -435
rect 1550 -1615 1560 -445
rect 1580 -1615 1590 -445
rect 1550 -1625 1590 -1615
rect 1650 -445 1690 -435
rect 1650 -1615 1660 -445
rect 1680 -1615 1690 -445
rect 1650 -1625 1690 -1615
rect 1750 -445 1790 -435
rect 1750 -1615 1760 -445
rect 1780 -1615 1790 -445
rect 1750 -1625 1790 -1615
rect 1850 -445 1990 -435
rect 1850 -1615 1860 -445
rect 1880 -1615 1910 -445
rect 1930 -1615 1960 -445
rect 1980 -1615 1990 -445
rect 1850 -1625 1990 -1615
rect 2050 -445 2090 -435
rect 2050 -1615 2060 -445
rect 2080 -1615 2090 -445
rect 2050 -1625 2090 -1615
rect 2150 -445 2190 -435
rect 2150 -1615 2160 -445
rect 2180 -1615 2190 -445
rect 2150 -1625 2190 -1615
rect 2250 -445 2290 -435
rect 2250 -1615 2260 -445
rect 2280 -1615 2290 -445
rect 2250 -1625 2290 -1615
rect 2350 -445 2390 -435
rect 2350 -1615 2360 -445
rect 2380 -1615 2390 -445
rect 2350 -1625 2390 -1615
rect 2450 -445 2490 -435
rect 2450 -1615 2460 -445
rect 2480 -1615 2490 -445
rect 2450 -1625 2490 -1615
rect 2530 -445 2620 -435
rect 2530 -1615 2540 -445
rect 2560 -1615 2590 -445
rect 2610 -1615 2620 -445
rect 2530 -1625 2620 -1615
rect 2680 -445 2720 -435
rect 2680 -1615 2690 -445
rect 2710 -1615 2720 -445
rect 2680 -1625 2720 -1615
rect 2760 -445 2850 -435
rect 2760 -1615 2770 -445
rect 2790 -1615 2820 -445
rect 2840 -1615 2850 -445
rect 2760 -1625 2850 -1615
rect 2910 -445 2950 -435
rect 2910 -1615 2920 -445
rect 2940 -1615 2950 -445
rect 2910 -1625 2950 -1615
rect 3015 -435 3035 -415
rect 3185 -390 3225 -380
rect 3185 -410 3195 -390
rect 3215 -410 3225 -390
rect 3185 -420 3225 -410
rect 3185 -435 3205 -420
rect 3015 -445 3055 -435
rect 3015 -1615 3025 -445
rect 3045 -1615 3055 -445
rect 3015 -1625 3055 -1615
rect 3115 -445 3205 -435
rect 3115 -1615 3125 -445
rect 3145 -1615 3175 -445
rect 3195 -1615 3205 -445
rect 3115 -1625 3205 -1615
rect 1250 -1675 1260 -1655
rect 1280 -1675 1290 -1655
rect 1250 -1685 1290 -1675
rect 1460 -1685 1480 -1625
rect 1660 -1685 1680 -1625
rect 2160 -1645 2180 -1625
rect 2540 -1645 2560 -1625
rect 2160 -1665 2560 -1645
rect 3115 -1655 3155 -1625
rect 3060 -1665 3155 -1655
rect 3060 -1685 3070 -1665
rect 1460 -1695 3070 -1685
rect 3100 -1675 3155 -1665
rect 3100 -1695 3110 -1675
rect 1460 -1705 3110 -1695
<< viali >>
rect 1245 -115 1265 1055
rect 1295 -115 1315 1055
rect 1795 -115 1815 1055
rect 1995 -115 2015 1055
rect 2045 -115 2065 1055
rect 2095 -115 2115 1055
rect 2495 -115 2515 1055
rect 2795 -115 2815 1055
rect 2845 -115 2865 1055
rect 3125 -115 3145 1055
rect 1260 -1615 1280 -445
rect 1360 -1615 1380 -445
rect 1860 -1615 1880 -445
rect 1910 -1615 1930 -445
rect 1960 -1615 1980 -445
rect 2460 -1615 2480 -445
rect 2770 -1615 2790 -445
rect 2820 -1615 2840 -445
<< metal1 >>
rect 1210 1055 3265 1065
rect 1210 -115 1245 1055
rect 1265 -115 1295 1055
rect 1315 -115 1795 1055
rect 1815 -115 1995 1055
rect 2015 -115 2045 1055
rect 2065 -115 2095 1055
rect 2115 -115 2495 1055
rect 2515 -115 2795 1055
rect 2815 -115 2845 1055
rect 2865 -115 3125 1055
rect 3145 -115 3265 1055
rect 1210 -125 3265 -115
rect 1210 -445 3265 -435
rect 1210 -1615 1260 -445
rect 1280 -1615 1360 -445
rect 1380 -1615 1860 -445
rect 1880 -1615 1910 -445
rect 1930 -1615 1960 -445
rect 1980 -1615 2460 -445
rect 2480 -1615 2770 -445
rect 2790 -1615 2820 -445
rect 2840 -1615 3265 -445
rect 1210 -1625 3265 -1615
<< labels >>
rlabel locali 1210 -155 1210 -155 7 Vb
rlabel metal1 1210 75 1210 75 7 VP
rlabel metal1 1210 -835 1210 -835 7 VN
rlabel locali 3265 -115 3265 -115 3 Vcp
rlabel locali 3265 -245 3265 -245 3 Vbn
rlabel locali 3265 -310 3265 -310 3 Vcn
<< end >>
