* SPICE3 file created from DFF.ext - technology: sky130A


* Top level circuit DFF

X0 a_n450_100# a_n500_n700# a_n470_n440# VN sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X1 VN Q Qn VN sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=9.5e+11p ps=5.9e+06u w=1e+06u l=150000u
X2 a_n40_380# Q Qn VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X3 Q Qn a_n40_380# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X4 Qn clk a_n500_n700# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1e+12p ps=6e+06u w=1e+06u l=600000u
X5 VP clk a_n40_380# VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_n450_100# a_n500_n700# VP VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_n470_n440# a_n450_100# a_n500_n700# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Q Qn VN VN sky130_fd_pr__nfet_01v8 ad=1e+12p pd=6e+06u as=0p ps=0u w=1e+06u l=150000u
X9 VP a_n450_100# a_n500_n700# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X10 Q clk a_n450_100# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=600000u
X11 a_n500_n700# clk Dn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5.5e+11p ps=3.1e+06u w=1e+06u l=600000u
X12 VN clk a_n470_n440# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 D clk a_n450_100# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=600000u
.end

